// Generator : SpinalHDL v1.8.0b    git head : 761a30e521263983ddf14de3592f7a9f38bf0589
// Component : MyTry
// Git hash  : 259ceaae35e16a989402949138e9eef49f0818f3

`timescale 1ns/1ps

module MyTry (
  input               io_a,
  output              io_b
);


  assign io_b = io_a;

endmodule
