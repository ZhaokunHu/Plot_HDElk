// Generator : SpinalHDL v1.8.0b    git head : 761a30e521263983ddf14de3592f7a9f38bf0589
// Component : top4
// Git hash  : c9998f03d07a31a5e92ff9ef47226a3ca5f7286c

`timescale 1ns/1ps

module top4 (
  input               io_a,
  output              io_b
);


  assign io_b = io_a;

endmodule
