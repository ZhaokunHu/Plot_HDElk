// Generator : SpinalHDL v1.8.0b    git head : 761a30e521263983ddf14de3592f7a9f38bf0589
// Component : TopLevel
// Git hash  : dc99cfcc67aa6033fefea7c05cf7cfef31e92939

`timescale 1ns/1ps

module TopLevel (
  input               KEY_Fn,
  input               CLK_50,
  input      [20:0]   COL,
  output     [5:0]    LED_A,
  output     [5:0]    ROW,
  output     [34:0]   LED_K,
  output              TXD,
  output              LED_R6,
  inout               PS2_CLK,
  inout               PS2_DAT,
  output              flash_dclk,
  output              flash_sce,
  output              flash_sdo,
  input               flash_data0
);
  localparam UartParityType_NONE = 2'd0;
  localparam UartParityType_EVEN = 2'd1;
  localparam UartParityType_ODD = 2'd2;
  localparam UartStopType_ONE = 1'd0;
  localparam UartStopType_TWO = 1'd1;

  wire                rstCtrl_io_externalReset;
  wire                core_reset_reset_n;
  wire                uartCtrl_2_io_read_ready;
  wire                clk50Area_hid_keyStatus_0_valid;
  wire                clk50Area_hid_keyStatus_0_payload;
  wire                clk50Area_hid_keyStatus_1_valid;
  wire                clk50Area_hid_keyStatus_1_payload;
  wire                clk50Area_hid_keyStatus_2_valid;
  wire                clk50Area_hid_keyStatus_2_payload;
  wire                clk50Area_hid_keyStatus_3_valid;
  wire                clk50Area_hid_keyStatus_3_payload;
  wire                clk50Area_hid_keyStatus_4_valid;
  wire                clk50Area_hid_keyStatus_4_payload;
  wire                clk50Area_hid_keyStatus_5_valid;
  wire                clk50Area_hid_keyStatus_5_payload;
  wire                clk50Area_hid_keyStatus_6_valid;
  wire                clk50Area_hid_keyStatus_6_payload;
  wire                clk50Area_hid_keyStatus_7_valid;
  wire                clk50Area_hid_keyStatus_7_payload;
  wire                clk50Area_hid_keyStatus_8_valid;
  wire                clk50Area_hid_keyStatus_8_payload;
  wire                clk50Area_hid_keyStatus_9_valid;
  wire                clk50Area_hid_keyStatus_9_payload;
  wire                clk50Area_hid_keyStatus_10_valid;
  wire                clk50Area_hid_keyStatus_10_payload;
  wire                clk50Area_hid_keyStatus_11_valid;
  wire                clk50Area_hid_keyStatus_11_payload;
  wire                clk50Area_hid_keyStatus_12_valid;
  wire                clk50Area_hid_keyStatus_12_payload;
  wire                clk50Area_hid_keyStatus_13_valid;
  wire                clk50Area_hid_keyStatus_13_payload;
  wire                clk50Area_hid_keyStatus_14_valid;
  wire                clk50Area_hid_keyStatus_14_payload;
  wire                clk50Area_hid_keyStatus_15_valid;
  wire                clk50Area_hid_keyStatus_15_payload;
  wire                clk50Area_hid_keyStatus_16_valid;
  wire                clk50Area_hid_keyStatus_16_payload;
  wire                clk50Area_hid_keyStatus_17_valid;
  wire                clk50Area_hid_keyStatus_17_payload;
  wire                clk50Area_hid_keyStatus_18_valid;
  wire                clk50Area_hid_keyStatus_18_payload;
  wire                clk50Area_hid_keyStatus_19_valid;
  wire                clk50Area_hid_keyStatus_19_payload;
  wire                clk50Area_hid_keyStatus_20_valid;
  wire                clk50Area_hid_keyStatus_20_payload;
  wire                clk50Area_hid_keyStatus_21_valid;
  wire                clk50Area_hid_keyStatus_21_payload;
  wire                clk50Area_hid_keyStatus_22_valid;
  wire                clk50Area_hid_keyStatus_22_payload;
  wire                clk50Area_hid_keyStatus_23_valid;
  wire                clk50Area_hid_keyStatus_23_payload;
  wire                clk50Area_hid_keyStatus_24_valid;
  wire                clk50Area_hid_keyStatus_24_payload;
  wire                clk50Area_hid_keyStatus_25_valid;
  wire                clk50Area_hid_keyStatus_25_payload;
  wire                clk50Area_hid_keyStatus_26_valid;
  wire                clk50Area_hid_keyStatus_26_payload;
  wire                clk50Area_hid_keyStatus_27_valid;
  wire                clk50Area_hid_keyStatus_27_payload;
  wire                clk50Area_hid_keyStatus_28_valid;
  wire                clk50Area_hid_keyStatus_28_payload;
  wire                clk50Area_hid_keyStatus_29_valid;
  wire                clk50Area_hid_keyStatus_29_payload;
  wire                clk50Area_hid_keyStatus_30_valid;
  wire                clk50Area_hid_keyStatus_30_payload;
  wire                clk50Area_hid_keyStatus_31_valid;
  wire                clk50Area_hid_keyStatus_31_payload;
  wire                clk50Area_hid_keyStatus_32_valid;
  wire                clk50Area_hid_keyStatus_32_payload;
  wire                clk50Area_hid_keyStatus_33_valid;
  wire                clk50Area_hid_keyStatus_33_payload;
  wire                clk50Area_hid_keyStatus_34_valid;
  wire                clk50Area_hid_keyStatus_34_payload;
  wire                clk50Area_hid_keyStatus_35_valid;
  wire                clk50Area_hid_keyStatus_35_payload;
  wire                clk50Area_hid_keyStatus_36_valid;
  wire                clk50Area_hid_keyStatus_36_payload;
  wire                clk50Area_hid_keyStatus_37_valid;
  wire                clk50Area_hid_keyStatus_37_payload;
  wire                clk50Area_hid_keyStatus_38_valid;
  wire                clk50Area_hid_keyStatus_38_payload;
  wire                clk50Area_hid_keyStatus_39_valid;
  wire                clk50Area_hid_keyStatus_39_payload;
  wire                clk50Area_hid_keyStatus_40_valid;
  wire                clk50Area_hid_keyStatus_40_payload;
  wire                clk50Area_hid_keyStatus_41_valid;
  wire                clk50Area_hid_keyStatus_41_payload;
  wire                clk50Area_hid_keyStatus_42_valid;
  wire                clk50Area_hid_keyStatus_42_payload;
  wire                clk50Area_hid_keyStatus_43_valid;
  wire                clk50Area_hid_keyStatus_43_payload;
  wire                clk50Area_hid_keyStatus_44_valid;
  wire                clk50Area_hid_keyStatus_44_payload;
  wire                clk50Area_hid_keyStatus_45_valid;
  wire                clk50Area_hid_keyStatus_45_payload;
  wire                clk50Area_hid_keyStatus_46_valid;
  wire                clk50Area_hid_keyStatus_46_payload;
  wire                clk50Area_hid_keyStatus_47_valid;
  wire                clk50Area_hid_keyStatus_47_payload;
  wire                clk50Area_hid_keyStatus_48_valid;
  wire                clk50Area_hid_keyStatus_48_payload;
  wire                clk50Area_hid_keyStatus_49_valid;
  wire                clk50Area_hid_keyStatus_49_payload;
  wire                clk50Area_hid_keyStatus_50_valid;
  wire                clk50Area_hid_keyStatus_50_payload;
  wire                clk50Area_hid_keyStatus_51_valid;
  wire                clk50Area_hid_keyStatus_51_payload;
  wire                clk50Area_hid_keyStatus_52_valid;
  wire                clk50Area_hid_keyStatus_52_payload;
  wire                clk50Area_hid_keyStatus_53_valid;
  wire                clk50Area_hid_keyStatus_53_payload;
  wire                clk50Area_hid_keyStatus_54_valid;
  wire                clk50Area_hid_keyStatus_54_payload;
  wire                clk50Area_hid_keyStatus_55_valid;
  wire                clk50Area_hid_keyStatus_55_payload;
  wire                clk50Area_hid_keyStatus_56_valid;
  wire                clk50Area_hid_keyStatus_56_payload;
  wire                clk50Area_hid_keyStatus_57_valid;
  wire                clk50Area_hid_keyStatus_57_payload;
  wire                clk50Area_hid_keyStatus_58_valid;
  wire                clk50Area_hid_keyStatus_58_payload;
  wire                clk50Area_hid_keyStatus_59_valid;
  wire                clk50Area_hid_keyStatus_59_payload;
  wire                clk50Area_hid_keyStatus_60_valid;
  wire                clk50Area_hid_keyStatus_60_payload;
  wire                clk50Area_hid_keyStatus_61_valid;
  wire                clk50Area_hid_keyStatus_61_payload;
  wire                clk50Area_hid_keyStatus_62_valid;
  wire                clk50Area_hid_keyStatus_62_payload;
  wire                clk50Area_hid_keyStatus_63_valid;
  wire                clk50Area_hid_keyStatus_63_payload;
  wire                clk50Area_hid_keyStatus_64_valid;
  wire                clk50Area_hid_keyStatus_64_payload;
  wire                clk50Area_hid_keyStatus_65_valid;
  wire                clk50Area_hid_keyStatus_65_payload;
  wire                clk50Area_hid_keyStatus_66_valid;
  wire                clk50Area_hid_keyStatus_66_payload;
  wire                clk50Area_hid_keyStatus_67_valid;
  wire                clk50Area_hid_keyStatus_67_payload;
  wire                clk50Area_hid_keyStatus_68_valid;
  wire                clk50Area_hid_keyStatus_68_payload;
  wire                clk50Area_hid_keyStatus_69_valid;
  wire                clk50Area_hid_keyStatus_69_payload;
  wire                clk50Area_hid_keyStatus_70_valid;
  wire                clk50Area_hid_keyStatus_70_payload;
  wire                clk50Area_hid_keyStatus_71_valid;
  wire                clk50Area_hid_keyStatus_71_payload;
  wire                clk50Area_hid_keyStatus_72_valid;
  wire                clk50Area_hid_keyStatus_72_payload;
  wire                clk50Area_hid_keyStatus_73_valid;
  wire                clk50Area_hid_keyStatus_73_payload;
  wire                clk50Area_hid_keyStatus_75_valid;
  wire                clk50Area_hid_keyStatus_75_payload;
  wire                clk50Area_hid_keyStatus_76_valid;
  wire                clk50Area_hid_keyStatus_76_payload;
  wire                clk50Area_hid_keyStatus_77_valid;
  wire                clk50Area_hid_keyStatus_77_payload;
  wire                clk50Area_hid_keyStatus_78_valid;
  wire                clk50Area_hid_keyStatus_78_payload;
  wire                clk50Area_hid_keyStatus_79_valid;
  wire                clk50Area_hid_keyStatus_79_payload;
  wire                clk50Area_hid_keyStatus_80_valid;
  wire                clk50Area_hid_keyStatus_80_payload;
  wire                clk50Area_hid_keyStatus_81_valid;
  wire                clk50Area_hid_keyStatus_81_payload;
  wire                clk50Area_hid_keyStatus_82_valid;
  wire                clk50Area_hid_keyStatus_82_payload;
  wire                clk50Area_hid_keyStatus_83_valid;
  wire                clk50Area_hid_keyStatus_83_payload;
  wire                clk50Area_hid_keyStatus_84_valid;
  wire                clk50Area_hid_keyStatus_84_payload;
  wire                clk50Area_hid_keyStatus_86_valid;
  wire                clk50Area_hid_keyStatus_86_payload;
  wire                clk50Area_hid_keyStatus_87_valid;
  wire                clk50Area_hid_keyStatus_87_payload;
  wire                clk50Area_hid_keyStatus_88_valid;
  wire                clk50Area_hid_keyStatus_88_payload;
  wire                clk50Area_hid_keyStatus_89_valid;
  wire                clk50Area_hid_keyStatus_89_payload;
  wire                clk50Area_hid_keyStatus_93_valid;
  wire                clk50Area_hid_keyStatus_93_payload;
  wire                clk50Area_hid_keyStatus_95_valid;
  wire                clk50Area_hid_keyStatus_95_payload;
  wire                clk50Area_hid_keyStatus_97_valid;
  wire                clk50Area_hid_keyStatus_97_payload;
  wire                clk50Area_hid_keyStatus_98_valid;
  wire                clk50Area_hid_keyStatus_98_payload;
  wire                clk50Area_hid_keyStatus_99_valid;
  wire                clk50Area_hid_keyStatus_99_payload;
  wire                clk50Area_hid_keyStatus_100_valid;
  wire                clk50Area_hid_keyStatus_100_payload;
  wire                clk50Area_hid_keyStatus_101_valid;
  wire                clk50Area_hid_keyStatus_101_payload;
  wire                clk50Area_hid_keyStatus_102_valid;
  wire                clk50Area_hid_keyStatus_102_payload;
  wire                pll100_c0;
  wire                pll100_locked;
  wire                rstCtrl_io_globalReset;
  wire                bufferCC_3_io_dataOut;
  wire                core_uart_txd;
  wire       [5:0]    core_io_row;
  wire       [34:0]   core_io_col;
  wire                core_flash_dclk;
  wire                core_flash_sce;
  wire                core_flash_sdo;
  wire       [5:0]    clk50Area_keyMatrix_ROW;
  wire                clk50Area_keyMatrix_scanIdx_valid;
  wire       [7:0]    clk50Area_keyMatrix_scanIdx_payload;
  wire                clk50Area_keyMatrix_keyStatus_0_valid;
  wire                clk50Area_keyMatrix_keyStatus_0_payload;
  wire                clk50Area_keyMatrix_keyStatus_1_valid;
  wire                clk50Area_keyMatrix_keyStatus_1_payload;
  wire                clk50Area_keyMatrix_keyStatus_2_valid;
  wire                clk50Area_keyMatrix_keyStatus_2_payload;
  wire                clk50Area_keyMatrix_keyStatus_3_valid;
  wire                clk50Area_keyMatrix_keyStatus_3_payload;
  wire                clk50Area_keyMatrix_keyStatus_4_valid;
  wire                clk50Area_keyMatrix_keyStatus_4_payload;
  wire                clk50Area_keyMatrix_keyStatus_5_valid;
  wire                clk50Area_keyMatrix_keyStatus_5_payload;
  wire                clk50Area_keyMatrix_keyStatus_6_valid;
  wire                clk50Area_keyMatrix_keyStatus_6_payload;
  wire                clk50Area_keyMatrix_keyStatus_7_valid;
  wire                clk50Area_keyMatrix_keyStatus_7_payload;
  wire                clk50Area_keyMatrix_keyStatus_8_valid;
  wire                clk50Area_keyMatrix_keyStatus_8_payload;
  wire                clk50Area_keyMatrix_keyStatus_9_valid;
  wire                clk50Area_keyMatrix_keyStatus_9_payload;
  wire                clk50Area_keyMatrix_keyStatus_10_valid;
  wire                clk50Area_keyMatrix_keyStatus_10_payload;
  wire                clk50Area_keyMatrix_keyStatus_11_valid;
  wire                clk50Area_keyMatrix_keyStatus_11_payload;
  wire                clk50Area_keyMatrix_keyStatus_12_valid;
  wire                clk50Area_keyMatrix_keyStatus_12_payload;
  wire                clk50Area_keyMatrix_keyStatus_13_valid;
  wire                clk50Area_keyMatrix_keyStatus_13_payload;
  wire                clk50Area_keyMatrix_keyStatus_14_valid;
  wire                clk50Area_keyMatrix_keyStatus_14_payload;
  wire                clk50Area_keyMatrix_keyStatus_15_valid;
  wire                clk50Area_keyMatrix_keyStatus_15_payload;
  wire                clk50Area_keyMatrix_keyStatus_16_valid;
  wire                clk50Area_keyMatrix_keyStatus_16_payload;
  wire                clk50Area_keyMatrix_keyStatus_17_valid;
  wire                clk50Area_keyMatrix_keyStatus_17_payload;
  wire                clk50Area_keyMatrix_keyStatus_18_valid;
  wire                clk50Area_keyMatrix_keyStatus_18_payload;
  wire                clk50Area_keyMatrix_keyStatus_19_valid;
  wire                clk50Area_keyMatrix_keyStatus_19_payload;
  wire                clk50Area_keyMatrix_keyStatus_20_valid;
  wire                clk50Area_keyMatrix_keyStatus_20_payload;
  wire                clk50Area_keyMatrix_keyStatus_21_valid;
  wire                clk50Area_keyMatrix_keyStatus_21_payload;
  wire                clk50Area_keyMatrix_keyStatus_22_valid;
  wire                clk50Area_keyMatrix_keyStatus_22_payload;
  wire                clk50Area_keyMatrix_keyStatus_23_valid;
  wire                clk50Area_keyMatrix_keyStatus_23_payload;
  wire                clk50Area_keyMatrix_keyStatus_24_valid;
  wire                clk50Area_keyMatrix_keyStatus_24_payload;
  wire                clk50Area_keyMatrix_keyStatus_25_valid;
  wire                clk50Area_keyMatrix_keyStatus_25_payload;
  wire                clk50Area_keyMatrix_keyStatus_26_valid;
  wire                clk50Area_keyMatrix_keyStatus_26_payload;
  wire                clk50Area_keyMatrix_keyStatus_27_valid;
  wire                clk50Area_keyMatrix_keyStatus_27_payload;
  wire                clk50Area_keyMatrix_keyStatus_28_valid;
  wire                clk50Area_keyMatrix_keyStatus_28_payload;
  wire                clk50Area_keyMatrix_keyStatus_29_valid;
  wire                clk50Area_keyMatrix_keyStatus_29_payload;
  wire                clk50Area_keyMatrix_keyStatus_30_valid;
  wire                clk50Area_keyMatrix_keyStatus_30_payload;
  wire                clk50Area_keyMatrix_keyStatus_31_valid;
  wire                clk50Area_keyMatrix_keyStatus_31_payload;
  wire                clk50Area_keyMatrix_keyStatus_32_valid;
  wire                clk50Area_keyMatrix_keyStatus_32_payload;
  wire                clk50Area_keyMatrix_keyStatus_33_valid;
  wire                clk50Area_keyMatrix_keyStatus_33_payload;
  wire                clk50Area_keyMatrix_keyStatus_34_valid;
  wire                clk50Area_keyMatrix_keyStatus_34_payload;
  wire                clk50Area_keyMatrix_keyStatus_35_valid;
  wire                clk50Area_keyMatrix_keyStatus_35_payload;
  wire                clk50Area_keyMatrix_keyStatus_36_valid;
  wire                clk50Area_keyMatrix_keyStatus_36_payload;
  wire                clk50Area_keyMatrix_keyStatus_37_valid;
  wire                clk50Area_keyMatrix_keyStatus_37_payload;
  wire                clk50Area_keyMatrix_keyStatus_38_valid;
  wire                clk50Area_keyMatrix_keyStatus_38_payload;
  wire                clk50Area_keyMatrix_keyStatus_39_valid;
  wire                clk50Area_keyMatrix_keyStatus_39_payload;
  wire                clk50Area_keyMatrix_keyStatus_40_valid;
  wire                clk50Area_keyMatrix_keyStatus_40_payload;
  wire                clk50Area_keyMatrix_keyStatus_41_valid;
  wire                clk50Area_keyMatrix_keyStatus_41_payload;
  wire                clk50Area_keyMatrix_keyStatus_42_valid;
  wire                clk50Area_keyMatrix_keyStatus_42_payload;
  wire                clk50Area_keyMatrix_keyStatus_43_valid;
  wire                clk50Area_keyMatrix_keyStatus_43_payload;
  wire                clk50Area_keyMatrix_keyStatus_44_valid;
  wire                clk50Area_keyMatrix_keyStatus_44_payload;
  wire                clk50Area_keyMatrix_keyStatus_45_valid;
  wire                clk50Area_keyMatrix_keyStatus_45_payload;
  wire                clk50Area_keyMatrix_keyStatus_46_valid;
  wire                clk50Area_keyMatrix_keyStatus_46_payload;
  wire                clk50Area_keyMatrix_keyStatus_47_valid;
  wire                clk50Area_keyMatrix_keyStatus_47_payload;
  wire                clk50Area_keyMatrix_keyStatus_48_valid;
  wire                clk50Area_keyMatrix_keyStatus_48_payload;
  wire                clk50Area_keyMatrix_keyStatus_49_valid;
  wire                clk50Area_keyMatrix_keyStatus_49_payload;
  wire                clk50Area_keyMatrix_keyStatus_50_valid;
  wire                clk50Area_keyMatrix_keyStatus_50_payload;
  wire                clk50Area_keyMatrix_keyStatus_51_valid;
  wire                clk50Area_keyMatrix_keyStatus_51_payload;
  wire                clk50Area_keyMatrix_keyStatus_52_valid;
  wire                clk50Area_keyMatrix_keyStatus_52_payload;
  wire                clk50Area_keyMatrix_keyStatus_53_valid;
  wire                clk50Area_keyMatrix_keyStatus_53_payload;
  wire                clk50Area_keyMatrix_keyStatus_54_valid;
  wire                clk50Area_keyMatrix_keyStatus_54_payload;
  wire                clk50Area_keyMatrix_keyStatus_55_valid;
  wire                clk50Area_keyMatrix_keyStatus_55_payload;
  wire                clk50Area_keyMatrix_keyStatus_56_valid;
  wire                clk50Area_keyMatrix_keyStatus_56_payload;
  wire                clk50Area_keyMatrix_keyStatus_57_valid;
  wire                clk50Area_keyMatrix_keyStatus_57_payload;
  wire                clk50Area_keyMatrix_keyStatus_58_valid;
  wire                clk50Area_keyMatrix_keyStatus_58_payload;
  wire                clk50Area_keyMatrix_keyStatus_59_valid;
  wire                clk50Area_keyMatrix_keyStatus_59_payload;
  wire                clk50Area_keyMatrix_keyStatus_60_valid;
  wire                clk50Area_keyMatrix_keyStatus_60_payload;
  wire                clk50Area_keyMatrix_keyStatus_61_valid;
  wire                clk50Area_keyMatrix_keyStatus_61_payload;
  wire                clk50Area_keyMatrix_keyStatus_62_valid;
  wire                clk50Area_keyMatrix_keyStatus_62_payload;
  wire                clk50Area_keyMatrix_keyStatus_63_valid;
  wire                clk50Area_keyMatrix_keyStatus_63_payload;
  wire                clk50Area_keyMatrix_keyStatus_64_valid;
  wire                clk50Area_keyMatrix_keyStatus_64_payload;
  wire                clk50Area_keyMatrix_keyStatus_65_valid;
  wire                clk50Area_keyMatrix_keyStatus_65_payload;
  wire                clk50Area_keyMatrix_keyStatus_66_valid;
  wire                clk50Area_keyMatrix_keyStatus_66_payload;
  wire                clk50Area_keyMatrix_keyStatus_67_valid;
  wire                clk50Area_keyMatrix_keyStatus_67_payload;
  wire                clk50Area_keyMatrix_keyStatus_68_valid;
  wire                clk50Area_keyMatrix_keyStatus_68_payload;
  wire                clk50Area_keyMatrix_keyStatus_69_valid;
  wire                clk50Area_keyMatrix_keyStatus_69_payload;
  wire                clk50Area_keyMatrix_keyStatus_70_valid;
  wire                clk50Area_keyMatrix_keyStatus_70_payload;
  wire                clk50Area_keyMatrix_keyStatus_71_valid;
  wire                clk50Area_keyMatrix_keyStatus_71_payload;
  wire                clk50Area_keyMatrix_keyStatus_72_valid;
  wire                clk50Area_keyMatrix_keyStatus_72_payload;
  wire                clk50Area_keyMatrix_keyStatus_73_valid;
  wire                clk50Area_keyMatrix_keyStatus_73_payload;
  wire                clk50Area_keyMatrix_keyStatus_74_valid;
  wire                clk50Area_keyMatrix_keyStatus_74_payload;
  wire                clk50Area_keyMatrix_keyStatus_75_valid;
  wire                clk50Area_keyMatrix_keyStatus_75_payload;
  wire                clk50Area_keyMatrix_keyStatus_76_valid;
  wire                clk50Area_keyMatrix_keyStatus_76_payload;
  wire                clk50Area_keyMatrix_keyStatus_77_valid;
  wire                clk50Area_keyMatrix_keyStatus_77_payload;
  wire                clk50Area_keyMatrix_keyStatus_78_valid;
  wire                clk50Area_keyMatrix_keyStatus_78_payload;
  wire                clk50Area_keyMatrix_keyStatus_79_valid;
  wire                clk50Area_keyMatrix_keyStatus_79_payload;
  wire                clk50Area_keyMatrix_keyStatus_80_valid;
  wire                clk50Area_keyMatrix_keyStatus_80_payload;
  wire                clk50Area_keyMatrix_keyStatus_81_valid;
  wire                clk50Area_keyMatrix_keyStatus_81_payload;
  wire                clk50Area_keyMatrix_keyStatus_82_valid;
  wire                clk50Area_keyMatrix_keyStatus_82_payload;
  wire                clk50Area_keyMatrix_keyStatus_83_valid;
  wire                clk50Area_keyMatrix_keyStatus_83_payload;
  wire                clk50Area_keyMatrix_keyStatus_84_valid;
  wire                clk50Area_keyMatrix_keyStatus_84_payload;
  wire                clk50Area_keyMatrix_keyStatus_85_valid;
  wire                clk50Area_keyMatrix_keyStatus_85_payload;
  wire                clk50Area_keyMatrix_keyStatus_86_valid;
  wire                clk50Area_keyMatrix_keyStatus_86_payload;
  wire                clk50Area_keyMatrix_keyStatus_87_valid;
  wire                clk50Area_keyMatrix_keyStatus_87_payload;
  wire                clk50Area_keyMatrix_keyStatus_88_valid;
  wire                clk50Area_keyMatrix_keyStatus_88_payload;
  wire                clk50Area_keyMatrix_keyStatus_89_valid;
  wire                clk50Area_keyMatrix_keyStatus_89_payload;
  wire                clk50Area_keyMatrix_keyStatus_90_valid;
  wire                clk50Area_keyMatrix_keyStatus_90_payload;
  wire                clk50Area_keyMatrix_keyStatus_91_valid;
  wire                clk50Area_keyMatrix_keyStatus_91_payload;
  wire                clk50Area_keyMatrix_keyStatus_92_valid;
  wire                clk50Area_keyMatrix_keyStatus_92_payload;
  wire                clk50Area_keyMatrix_keyStatus_93_valid;
  wire                clk50Area_keyMatrix_keyStatus_93_payload;
  wire                clk50Area_keyMatrix_keyStatus_94_valid;
  wire                clk50Area_keyMatrix_keyStatus_94_payload;
  wire                clk50Area_keyMatrix_keyStatus_95_valid;
  wire                clk50Area_keyMatrix_keyStatus_95_payload;
  wire                clk50Area_keyMatrix_keyStatus_96_valid;
  wire                clk50Area_keyMatrix_keyStatus_96_payload;
  wire                clk50Area_keyMatrix_keyStatus_97_valid;
  wire                clk50Area_keyMatrix_keyStatus_97_payload;
  wire                clk50Area_keyMatrix_keyStatus_98_valid;
  wire                clk50Area_keyMatrix_keyStatus_98_payload;
  wire                clk50Area_keyMatrix_keyStatus_99_valid;
  wire                clk50Area_keyMatrix_keyStatus_99_payload;
  wire                clk50Area_keyMatrix_keyStatus_100_valid;
  wire                clk50Area_keyMatrix_keyStatus_100_payload;
  wire                clk50Area_keyMatrix_keyStatus_101_valid;
  wire                clk50Area_keyMatrix_keyStatus_101_payload;
  wire                clk50Area_keyMatrix_keyStatus_102_valid;
  wire                clk50Area_keyMatrix_keyStatus_102_payload;
  wire                uartCtrl_2_io_write_ready;
  wire                uartCtrl_2_io_read_valid;
  wire       [7:0]    uartCtrl_2_io_read_payload;
  wire                uartCtrl_2_io_uart_txd;
  wire                uartCtrl_2_io_readError;
  wire                uartCtrl_2_io_readBreak;
  wire                clk50Area_hid_TXD;
  reg                 _zz_LED_R6;
  wire                _zz_1;
  reg        [7:0]    toplevel_clk50Area_keyMatrix_scanIdx_payload_regNextWhen;
  reg                 _zz_io_write_valid;

  pll pll100 (
    .inclk0 (CLK_50       ), //i
    .c0     (pll100_c0    ), //o
    .locked (pll100_locked)  //o
  );
  ResetController rstCtrl (
    .io_clock         (CLK_50                  ), //i
    .io_externalReset (rstCtrl_io_externalReset), //i
    .io_globalReset   (rstCtrl_io_globalReset  )  //o
  );
  BufferCC bufferCC_3 (
    .io_dataIn  (1'b0                 ), //i
    .io_dataOut (bufferCC_3_io_dataOut), //o
    .CLK_50     (CLK_50               ), //i
    ._zz_1      (_zz_1                )  //i
  );
  kbd104 core (
    .clk_clk       (pll100_c0             ), //i
    .reset_reset_n (core_reset_reset_n    ), //i
    .uart_txd      (core_uart_txd         ), //o
    .uart_rxd      (uartCtrl_2_io_uart_txd), //i
    .io_row        (core_io_row[5:0]      ), //o
    .io_col        (core_io_col[34:0]     ), //o
    .flash_dclk    (core_flash_dclk       ), //o
    .flash_sce     (core_flash_sce        ), //o
    .flash_sdo     (core_flash_sdo        ), //o
    .flash_data0   (flash_data0           )  //i
  );
  KeyMatrix clk50Area_keyMatrix (
    .enabled               (1'b1                                     ), //i
    .COL                   (COL[20:0]                                ), //i
    .ROW                   (clk50Area_keyMatrix_ROW[5:0]             ), //o
    .scanIdx_valid         (clk50Area_keyMatrix_scanIdx_valid        ), //o
    .scanIdx_payload       (clk50Area_keyMatrix_scanIdx_payload[7:0] ), //o
    .keyStatus_0_valid     (clk50Area_keyMatrix_keyStatus_0_valid    ), //o
    .keyStatus_0_payload   (clk50Area_keyMatrix_keyStatus_0_payload  ), //o
    .keyStatus_1_valid     (clk50Area_keyMatrix_keyStatus_1_valid    ), //o
    .keyStatus_1_payload   (clk50Area_keyMatrix_keyStatus_1_payload  ), //o
    .keyStatus_2_valid     (clk50Area_keyMatrix_keyStatus_2_valid    ), //o
    .keyStatus_2_payload   (clk50Area_keyMatrix_keyStatus_2_payload  ), //o
    .keyStatus_3_valid     (clk50Area_keyMatrix_keyStatus_3_valid    ), //o
    .keyStatus_3_payload   (clk50Area_keyMatrix_keyStatus_3_payload  ), //o
    .keyStatus_4_valid     (clk50Area_keyMatrix_keyStatus_4_valid    ), //o
    .keyStatus_4_payload   (clk50Area_keyMatrix_keyStatus_4_payload  ), //o
    .keyStatus_5_valid     (clk50Area_keyMatrix_keyStatus_5_valid    ), //o
    .keyStatus_5_payload   (clk50Area_keyMatrix_keyStatus_5_payload  ), //o
    .keyStatus_6_valid     (clk50Area_keyMatrix_keyStatus_6_valid    ), //o
    .keyStatus_6_payload   (clk50Area_keyMatrix_keyStatus_6_payload  ), //o
    .keyStatus_7_valid     (clk50Area_keyMatrix_keyStatus_7_valid    ), //o
    .keyStatus_7_payload   (clk50Area_keyMatrix_keyStatus_7_payload  ), //o
    .keyStatus_8_valid     (clk50Area_keyMatrix_keyStatus_8_valid    ), //o
    .keyStatus_8_payload   (clk50Area_keyMatrix_keyStatus_8_payload  ), //o
    .keyStatus_9_valid     (clk50Area_keyMatrix_keyStatus_9_valid    ), //o
    .keyStatus_9_payload   (clk50Area_keyMatrix_keyStatus_9_payload  ), //o
    .keyStatus_10_valid    (clk50Area_keyMatrix_keyStatus_10_valid   ), //o
    .keyStatus_10_payload  (clk50Area_keyMatrix_keyStatus_10_payload ), //o
    .keyStatus_11_valid    (clk50Area_keyMatrix_keyStatus_11_valid   ), //o
    .keyStatus_11_payload  (clk50Area_keyMatrix_keyStatus_11_payload ), //o
    .keyStatus_12_valid    (clk50Area_keyMatrix_keyStatus_12_valid   ), //o
    .keyStatus_12_payload  (clk50Area_keyMatrix_keyStatus_12_payload ), //o
    .keyStatus_13_valid    (clk50Area_keyMatrix_keyStatus_13_valid   ), //o
    .keyStatus_13_payload  (clk50Area_keyMatrix_keyStatus_13_payload ), //o
    .keyStatus_14_valid    (clk50Area_keyMatrix_keyStatus_14_valid   ), //o
    .keyStatus_14_payload  (clk50Area_keyMatrix_keyStatus_14_payload ), //o
    .keyStatus_15_valid    (clk50Area_keyMatrix_keyStatus_15_valid   ), //o
    .keyStatus_15_payload  (clk50Area_keyMatrix_keyStatus_15_payload ), //o
    .keyStatus_16_valid    (clk50Area_keyMatrix_keyStatus_16_valid   ), //o
    .keyStatus_16_payload  (clk50Area_keyMatrix_keyStatus_16_payload ), //o
    .keyStatus_17_valid    (clk50Area_keyMatrix_keyStatus_17_valid   ), //o
    .keyStatus_17_payload  (clk50Area_keyMatrix_keyStatus_17_payload ), //o
    .keyStatus_18_valid    (clk50Area_keyMatrix_keyStatus_18_valid   ), //o
    .keyStatus_18_payload  (clk50Area_keyMatrix_keyStatus_18_payload ), //o
    .keyStatus_19_valid    (clk50Area_keyMatrix_keyStatus_19_valid   ), //o
    .keyStatus_19_payload  (clk50Area_keyMatrix_keyStatus_19_payload ), //o
    .keyStatus_20_valid    (clk50Area_keyMatrix_keyStatus_20_valid   ), //o
    .keyStatus_20_payload  (clk50Area_keyMatrix_keyStatus_20_payload ), //o
    .keyStatus_21_valid    (clk50Area_keyMatrix_keyStatus_21_valid   ), //o
    .keyStatus_21_payload  (clk50Area_keyMatrix_keyStatus_21_payload ), //o
    .keyStatus_22_valid    (clk50Area_keyMatrix_keyStatus_22_valid   ), //o
    .keyStatus_22_payload  (clk50Area_keyMatrix_keyStatus_22_payload ), //o
    .keyStatus_23_valid    (clk50Area_keyMatrix_keyStatus_23_valid   ), //o
    .keyStatus_23_payload  (clk50Area_keyMatrix_keyStatus_23_payload ), //o
    .keyStatus_24_valid    (clk50Area_keyMatrix_keyStatus_24_valid   ), //o
    .keyStatus_24_payload  (clk50Area_keyMatrix_keyStatus_24_payload ), //o
    .keyStatus_25_valid    (clk50Area_keyMatrix_keyStatus_25_valid   ), //o
    .keyStatus_25_payload  (clk50Area_keyMatrix_keyStatus_25_payload ), //o
    .keyStatus_26_valid    (clk50Area_keyMatrix_keyStatus_26_valid   ), //o
    .keyStatus_26_payload  (clk50Area_keyMatrix_keyStatus_26_payload ), //o
    .keyStatus_27_valid    (clk50Area_keyMatrix_keyStatus_27_valid   ), //o
    .keyStatus_27_payload  (clk50Area_keyMatrix_keyStatus_27_payload ), //o
    .keyStatus_28_valid    (clk50Area_keyMatrix_keyStatus_28_valid   ), //o
    .keyStatus_28_payload  (clk50Area_keyMatrix_keyStatus_28_payload ), //o
    .keyStatus_29_valid    (clk50Area_keyMatrix_keyStatus_29_valid   ), //o
    .keyStatus_29_payload  (clk50Area_keyMatrix_keyStatus_29_payload ), //o
    .keyStatus_30_valid    (clk50Area_keyMatrix_keyStatus_30_valid   ), //o
    .keyStatus_30_payload  (clk50Area_keyMatrix_keyStatus_30_payload ), //o
    .keyStatus_31_valid    (clk50Area_keyMatrix_keyStatus_31_valid   ), //o
    .keyStatus_31_payload  (clk50Area_keyMatrix_keyStatus_31_payload ), //o
    .keyStatus_32_valid    (clk50Area_keyMatrix_keyStatus_32_valid   ), //o
    .keyStatus_32_payload  (clk50Area_keyMatrix_keyStatus_32_payload ), //o
    .keyStatus_33_valid    (clk50Area_keyMatrix_keyStatus_33_valid   ), //o
    .keyStatus_33_payload  (clk50Area_keyMatrix_keyStatus_33_payload ), //o
    .keyStatus_34_valid    (clk50Area_keyMatrix_keyStatus_34_valid   ), //o
    .keyStatus_34_payload  (clk50Area_keyMatrix_keyStatus_34_payload ), //o
    .keyStatus_35_valid    (clk50Area_keyMatrix_keyStatus_35_valid   ), //o
    .keyStatus_35_payload  (clk50Area_keyMatrix_keyStatus_35_payload ), //o
    .keyStatus_36_valid    (clk50Area_keyMatrix_keyStatus_36_valid   ), //o
    .keyStatus_36_payload  (clk50Area_keyMatrix_keyStatus_36_payload ), //o
    .keyStatus_37_valid    (clk50Area_keyMatrix_keyStatus_37_valid   ), //o
    .keyStatus_37_payload  (clk50Area_keyMatrix_keyStatus_37_payload ), //o
    .keyStatus_38_valid    (clk50Area_keyMatrix_keyStatus_38_valid   ), //o
    .keyStatus_38_payload  (clk50Area_keyMatrix_keyStatus_38_payload ), //o
    .keyStatus_39_valid    (clk50Area_keyMatrix_keyStatus_39_valid   ), //o
    .keyStatus_39_payload  (clk50Area_keyMatrix_keyStatus_39_payload ), //o
    .keyStatus_40_valid    (clk50Area_keyMatrix_keyStatus_40_valid   ), //o
    .keyStatus_40_payload  (clk50Area_keyMatrix_keyStatus_40_payload ), //o
    .keyStatus_41_valid    (clk50Area_keyMatrix_keyStatus_41_valid   ), //o
    .keyStatus_41_payload  (clk50Area_keyMatrix_keyStatus_41_payload ), //o
    .keyStatus_42_valid    (clk50Area_keyMatrix_keyStatus_42_valid   ), //o
    .keyStatus_42_payload  (clk50Area_keyMatrix_keyStatus_42_payload ), //o
    .keyStatus_43_valid    (clk50Area_keyMatrix_keyStatus_43_valid   ), //o
    .keyStatus_43_payload  (clk50Area_keyMatrix_keyStatus_43_payload ), //o
    .keyStatus_44_valid    (clk50Area_keyMatrix_keyStatus_44_valid   ), //o
    .keyStatus_44_payload  (clk50Area_keyMatrix_keyStatus_44_payload ), //o
    .keyStatus_45_valid    (clk50Area_keyMatrix_keyStatus_45_valid   ), //o
    .keyStatus_45_payload  (clk50Area_keyMatrix_keyStatus_45_payload ), //o
    .keyStatus_46_valid    (clk50Area_keyMatrix_keyStatus_46_valid   ), //o
    .keyStatus_46_payload  (clk50Area_keyMatrix_keyStatus_46_payload ), //o
    .keyStatus_47_valid    (clk50Area_keyMatrix_keyStatus_47_valid   ), //o
    .keyStatus_47_payload  (clk50Area_keyMatrix_keyStatus_47_payload ), //o
    .keyStatus_48_valid    (clk50Area_keyMatrix_keyStatus_48_valid   ), //o
    .keyStatus_48_payload  (clk50Area_keyMatrix_keyStatus_48_payload ), //o
    .keyStatus_49_valid    (clk50Area_keyMatrix_keyStatus_49_valid   ), //o
    .keyStatus_49_payload  (clk50Area_keyMatrix_keyStatus_49_payload ), //o
    .keyStatus_50_valid    (clk50Area_keyMatrix_keyStatus_50_valid   ), //o
    .keyStatus_50_payload  (clk50Area_keyMatrix_keyStatus_50_payload ), //o
    .keyStatus_51_valid    (clk50Area_keyMatrix_keyStatus_51_valid   ), //o
    .keyStatus_51_payload  (clk50Area_keyMatrix_keyStatus_51_payload ), //o
    .keyStatus_52_valid    (clk50Area_keyMatrix_keyStatus_52_valid   ), //o
    .keyStatus_52_payload  (clk50Area_keyMatrix_keyStatus_52_payload ), //o
    .keyStatus_53_valid    (clk50Area_keyMatrix_keyStatus_53_valid   ), //o
    .keyStatus_53_payload  (clk50Area_keyMatrix_keyStatus_53_payload ), //o
    .keyStatus_54_valid    (clk50Area_keyMatrix_keyStatus_54_valid   ), //o
    .keyStatus_54_payload  (clk50Area_keyMatrix_keyStatus_54_payload ), //o
    .keyStatus_55_valid    (clk50Area_keyMatrix_keyStatus_55_valid   ), //o
    .keyStatus_55_payload  (clk50Area_keyMatrix_keyStatus_55_payload ), //o
    .keyStatus_56_valid    (clk50Area_keyMatrix_keyStatus_56_valid   ), //o
    .keyStatus_56_payload  (clk50Area_keyMatrix_keyStatus_56_payload ), //o
    .keyStatus_57_valid    (clk50Area_keyMatrix_keyStatus_57_valid   ), //o
    .keyStatus_57_payload  (clk50Area_keyMatrix_keyStatus_57_payload ), //o
    .keyStatus_58_valid    (clk50Area_keyMatrix_keyStatus_58_valid   ), //o
    .keyStatus_58_payload  (clk50Area_keyMatrix_keyStatus_58_payload ), //o
    .keyStatus_59_valid    (clk50Area_keyMatrix_keyStatus_59_valid   ), //o
    .keyStatus_59_payload  (clk50Area_keyMatrix_keyStatus_59_payload ), //o
    .keyStatus_60_valid    (clk50Area_keyMatrix_keyStatus_60_valid   ), //o
    .keyStatus_60_payload  (clk50Area_keyMatrix_keyStatus_60_payload ), //o
    .keyStatus_61_valid    (clk50Area_keyMatrix_keyStatus_61_valid   ), //o
    .keyStatus_61_payload  (clk50Area_keyMatrix_keyStatus_61_payload ), //o
    .keyStatus_62_valid    (clk50Area_keyMatrix_keyStatus_62_valid   ), //o
    .keyStatus_62_payload  (clk50Area_keyMatrix_keyStatus_62_payload ), //o
    .keyStatus_63_valid    (clk50Area_keyMatrix_keyStatus_63_valid   ), //o
    .keyStatus_63_payload  (clk50Area_keyMatrix_keyStatus_63_payload ), //o
    .keyStatus_64_valid    (clk50Area_keyMatrix_keyStatus_64_valid   ), //o
    .keyStatus_64_payload  (clk50Area_keyMatrix_keyStatus_64_payload ), //o
    .keyStatus_65_valid    (clk50Area_keyMatrix_keyStatus_65_valid   ), //o
    .keyStatus_65_payload  (clk50Area_keyMatrix_keyStatus_65_payload ), //o
    .keyStatus_66_valid    (clk50Area_keyMatrix_keyStatus_66_valid   ), //o
    .keyStatus_66_payload  (clk50Area_keyMatrix_keyStatus_66_payload ), //o
    .keyStatus_67_valid    (clk50Area_keyMatrix_keyStatus_67_valid   ), //o
    .keyStatus_67_payload  (clk50Area_keyMatrix_keyStatus_67_payload ), //o
    .keyStatus_68_valid    (clk50Area_keyMatrix_keyStatus_68_valid   ), //o
    .keyStatus_68_payload  (clk50Area_keyMatrix_keyStatus_68_payload ), //o
    .keyStatus_69_valid    (clk50Area_keyMatrix_keyStatus_69_valid   ), //o
    .keyStatus_69_payload  (clk50Area_keyMatrix_keyStatus_69_payload ), //o
    .keyStatus_70_valid    (clk50Area_keyMatrix_keyStatus_70_valid   ), //o
    .keyStatus_70_payload  (clk50Area_keyMatrix_keyStatus_70_payload ), //o
    .keyStatus_71_valid    (clk50Area_keyMatrix_keyStatus_71_valid   ), //o
    .keyStatus_71_payload  (clk50Area_keyMatrix_keyStatus_71_payload ), //o
    .keyStatus_72_valid    (clk50Area_keyMatrix_keyStatus_72_valid   ), //o
    .keyStatus_72_payload  (clk50Area_keyMatrix_keyStatus_72_payload ), //o
    .keyStatus_73_valid    (clk50Area_keyMatrix_keyStatus_73_valid   ), //o
    .keyStatus_73_payload  (clk50Area_keyMatrix_keyStatus_73_payload ), //o
    .keyStatus_74_valid    (clk50Area_keyMatrix_keyStatus_74_valid   ), //o
    .keyStatus_74_payload  (clk50Area_keyMatrix_keyStatus_74_payload ), //o
    .keyStatus_75_valid    (clk50Area_keyMatrix_keyStatus_75_valid   ), //o
    .keyStatus_75_payload  (clk50Area_keyMatrix_keyStatus_75_payload ), //o
    .keyStatus_76_valid    (clk50Area_keyMatrix_keyStatus_76_valid   ), //o
    .keyStatus_76_payload  (clk50Area_keyMatrix_keyStatus_76_payload ), //o
    .keyStatus_77_valid    (clk50Area_keyMatrix_keyStatus_77_valid   ), //o
    .keyStatus_77_payload  (clk50Area_keyMatrix_keyStatus_77_payload ), //o
    .keyStatus_78_valid    (clk50Area_keyMatrix_keyStatus_78_valid   ), //o
    .keyStatus_78_payload  (clk50Area_keyMatrix_keyStatus_78_payload ), //o
    .keyStatus_79_valid    (clk50Area_keyMatrix_keyStatus_79_valid   ), //o
    .keyStatus_79_payload  (clk50Area_keyMatrix_keyStatus_79_payload ), //o
    .keyStatus_80_valid    (clk50Area_keyMatrix_keyStatus_80_valid   ), //o
    .keyStatus_80_payload  (clk50Area_keyMatrix_keyStatus_80_payload ), //o
    .keyStatus_81_valid    (clk50Area_keyMatrix_keyStatus_81_valid   ), //o
    .keyStatus_81_payload  (clk50Area_keyMatrix_keyStatus_81_payload ), //o
    .keyStatus_82_valid    (clk50Area_keyMatrix_keyStatus_82_valid   ), //o
    .keyStatus_82_payload  (clk50Area_keyMatrix_keyStatus_82_payload ), //o
    .keyStatus_83_valid    (clk50Area_keyMatrix_keyStatus_83_valid   ), //o
    .keyStatus_83_payload  (clk50Area_keyMatrix_keyStatus_83_payload ), //o
    .keyStatus_84_valid    (clk50Area_keyMatrix_keyStatus_84_valid   ), //o
    .keyStatus_84_payload  (clk50Area_keyMatrix_keyStatus_84_payload ), //o
    .keyStatus_85_valid    (clk50Area_keyMatrix_keyStatus_85_valid   ), //o
    .keyStatus_85_payload  (clk50Area_keyMatrix_keyStatus_85_payload ), //o
    .keyStatus_86_valid    (clk50Area_keyMatrix_keyStatus_86_valid   ), //o
    .keyStatus_86_payload  (clk50Area_keyMatrix_keyStatus_86_payload ), //o
    .keyStatus_87_valid    (clk50Area_keyMatrix_keyStatus_87_valid   ), //o
    .keyStatus_87_payload  (clk50Area_keyMatrix_keyStatus_87_payload ), //o
    .keyStatus_88_valid    (clk50Area_keyMatrix_keyStatus_88_valid   ), //o
    .keyStatus_88_payload  (clk50Area_keyMatrix_keyStatus_88_payload ), //o
    .keyStatus_89_valid    (clk50Area_keyMatrix_keyStatus_89_valid   ), //o
    .keyStatus_89_payload  (clk50Area_keyMatrix_keyStatus_89_payload ), //o
    .keyStatus_90_valid    (clk50Area_keyMatrix_keyStatus_90_valid   ), //o
    .keyStatus_90_payload  (clk50Area_keyMatrix_keyStatus_90_payload ), //o
    .keyStatus_91_valid    (clk50Area_keyMatrix_keyStatus_91_valid   ), //o
    .keyStatus_91_payload  (clk50Area_keyMatrix_keyStatus_91_payload ), //o
    .keyStatus_92_valid    (clk50Area_keyMatrix_keyStatus_92_valid   ), //o
    .keyStatus_92_payload  (clk50Area_keyMatrix_keyStatus_92_payload ), //o
    .keyStatus_93_valid    (clk50Area_keyMatrix_keyStatus_93_valid   ), //o
    .keyStatus_93_payload  (clk50Area_keyMatrix_keyStatus_93_payload ), //o
    .keyStatus_94_valid    (clk50Area_keyMatrix_keyStatus_94_valid   ), //o
    .keyStatus_94_payload  (clk50Area_keyMatrix_keyStatus_94_payload ), //o
    .keyStatus_95_valid    (clk50Area_keyMatrix_keyStatus_95_valid   ), //o
    .keyStatus_95_payload  (clk50Area_keyMatrix_keyStatus_95_payload ), //o
    .keyStatus_96_valid    (clk50Area_keyMatrix_keyStatus_96_valid   ), //o
    .keyStatus_96_payload  (clk50Area_keyMatrix_keyStatus_96_payload ), //o
    .keyStatus_97_valid    (clk50Area_keyMatrix_keyStatus_97_valid   ), //o
    .keyStatus_97_payload  (clk50Area_keyMatrix_keyStatus_97_payload ), //o
    .keyStatus_98_valid    (clk50Area_keyMatrix_keyStatus_98_valid   ), //o
    .keyStatus_98_payload  (clk50Area_keyMatrix_keyStatus_98_payload ), //o
    .keyStatus_99_valid    (clk50Area_keyMatrix_keyStatus_99_valid   ), //o
    .keyStatus_99_payload  (clk50Area_keyMatrix_keyStatus_99_payload ), //o
    .keyStatus_100_valid   (clk50Area_keyMatrix_keyStatus_100_valid  ), //o
    .keyStatus_100_payload (clk50Area_keyMatrix_keyStatus_100_payload), //o
    .keyStatus_101_valid   (clk50Area_keyMatrix_keyStatus_101_valid  ), //o
    .keyStatus_101_payload (clk50Area_keyMatrix_keyStatus_101_payload), //o
    .keyStatus_102_valid   (clk50Area_keyMatrix_keyStatus_102_valid  ), //o
    .keyStatus_102_payload (clk50Area_keyMatrix_keyStatus_102_payload), //o
    ._zz_LED_R6            (_zz_LED_R6                               ), //i
    .CLK_50                (CLK_50                                   )  //i
  );
  UartCtrl_1 uartCtrl_2 (
    .io_config_frame_dataLength (3'b111                                                       ), //i
    .io_config_frame_stop       (UartStopType_ONE                                             ), //i
    .io_config_frame_parity     (UartParityType_NONE                                          ), //i
    .io_config_clockDivider     (20'h00035                                                    ), //i
    .io_write_valid             (_zz_io_write_valid                                           ), //i
    .io_write_ready             (uartCtrl_2_io_write_ready                                    ), //o
    .io_write_payload           (toplevel_clk50Area_keyMatrix_scanIdx_payload_regNextWhen[7:0]), //i
    .io_read_valid              (uartCtrl_2_io_read_valid                                     ), //o
    .io_read_ready              (uartCtrl_2_io_read_ready                                     ), //i
    .io_read_payload            (uartCtrl_2_io_read_payload[7:0]                              ), //o
    .io_uart_txd                (uartCtrl_2_io_uart_txd                                       ), //o
    .io_uart_rxd                (1'b1                                                         ), //i
    .io_readError               (uartCtrl_2_io_readError                                      ), //o
    .io_writeBreak              (1'b0                                                         ), //i
    .io_readBreak               (uartCtrl_2_io_readBreak                                      ), //o
    .CLK_50                     (CLK_50                                                       ), //i
    ._zz_LED_R6                 (_zz_LED_R6                                                   )  //i
  );
  HID clk50Area_hid (
    .TXD                   (clk50Area_hid_TXD                       ), //o
    .scanIdx_valid         (clk50Area_keyMatrix_scanIdx_valid       ), //i
    .scanIdx_payload       (clk50Area_keyMatrix_scanIdx_payload[7:0]), //i
    .keyStatus_0_valid     (clk50Area_hid_keyStatus_0_valid         ), //i
    .keyStatus_0_payload   (clk50Area_hid_keyStatus_0_payload       ), //i
    .keyStatus_1_valid     (clk50Area_hid_keyStatus_1_valid         ), //i
    .keyStatus_1_payload   (clk50Area_hid_keyStatus_1_payload       ), //i
    .keyStatus_2_valid     (clk50Area_hid_keyStatus_2_valid         ), //i
    .keyStatus_2_payload   (clk50Area_hid_keyStatus_2_payload       ), //i
    .keyStatus_3_valid     (clk50Area_hid_keyStatus_3_valid         ), //i
    .keyStatus_3_payload   (clk50Area_hid_keyStatus_3_payload       ), //i
    .keyStatus_4_valid     (clk50Area_hid_keyStatus_4_valid         ), //i
    .keyStatus_4_payload   (clk50Area_hid_keyStatus_4_payload       ), //i
    .keyStatus_5_valid     (clk50Area_hid_keyStatus_5_valid         ), //i
    .keyStatus_5_payload   (clk50Area_hid_keyStatus_5_payload       ), //i
    .keyStatus_6_valid     (clk50Area_hid_keyStatus_6_valid         ), //i
    .keyStatus_6_payload   (clk50Area_hid_keyStatus_6_payload       ), //i
    .keyStatus_7_valid     (clk50Area_hid_keyStatus_7_valid         ), //i
    .keyStatus_7_payload   (clk50Area_hid_keyStatus_7_payload       ), //i
    .keyStatus_8_valid     (clk50Area_hid_keyStatus_8_valid         ), //i
    .keyStatus_8_payload   (clk50Area_hid_keyStatus_8_payload       ), //i
    .keyStatus_9_valid     (clk50Area_hid_keyStatus_9_valid         ), //i
    .keyStatus_9_payload   (clk50Area_hid_keyStatus_9_payload       ), //i
    .keyStatus_10_valid    (clk50Area_hid_keyStatus_10_valid        ), //i
    .keyStatus_10_payload  (clk50Area_hid_keyStatus_10_payload      ), //i
    .keyStatus_11_valid    (clk50Area_hid_keyStatus_11_valid        ), //i
    .keyStatus_11_payload  (clk50Area_hid_keyStatus_11_payload      ), //i
    .keyStatus_12_valid    (clk50Area_hid_keyStatus_12_valid        ), //i
    .keyStatus_12_payload  (clk50Area_hid_keyStatus_12_payload      ), //i
    .keyStatus_13_valid    (clk50Area_hid_keyStatus_13_valid        ), //i
    .keyStatus_13_payload  (clk50Area_hid_keyStatus_13_payload      ), //i
    .keyStatus_14_valid    (clk50Area_hid_keyStatus_14_valid        ), //i
    .keyStatus_14_payload  (clk50Area_hid_keyStatus_14_payload      ), //i
    .keyStatus_15_valid    (clk50Area_hid_keyStatus_15_valid        ), //i
    .keyStatus_15_payload  (clk50Area_hid_keyStatus_15_payload      ), //i
    .keyStatus_16_valid    (clk50Area_hid_keyStatus_16_valid        ), //i
    .keyStatus_16_payload  (clk50Area_hid_keyStatus_16_payload      ), //i
    .keyStatus_17_valid    (clk50Area_hid_keyStatus_17_valid        ), //i
    .keyStatus_17_payload  (clk50Area_hid_keyStatus_17_payload      ), //i
    .keyStatus_18_valid    (clk50Area_hid_keyStatus_18_valid        ), //i
    .keyStatus_18_payload  (clk50Area_hid_keyStatus_18_payload      ), //i
    .keyStatus_19_valid    (clk50Area_hid_keyStatus_19_valid        ), //i
    .keyStatus_19_payload  (clk50Area_hid_keyStatus_19_payload      ), //i
    .keyStatus_20_valid    (clk50Area_hid_keyStatus_20_valid        ), //i
    .keyStatus_20_payload  (clk50Area_hid_keyStatus_20_payload      ), //i
    .keyStatus_21_valid    (clk50Area_hid_keyStatus_21_valid        ), //i
    .keyStatus_21_payload  (clk50Area_hid_keyStatus_21_payload      ), //i
    .keyStatus_22_valid    (clk50Area_hid_keyStatus_22_valid        ), //i
    .keyStatus_22_payload  (clk50Area_hid_keyStatus_22_payload      ), //i
    .keyStatus_23_valid    (clk50Area_hid_keyStatus_23_valid        ), //i
    .keyStatus_23_payload  (clk50Area_hid_keyStatus_23_payload      ), //i
    .keyStatus_24_valid    (clk50Area_hid_keyStatus_24_valid        ), //i
    .keyStatus_24_payload  (clk50Area_hid_keyStatus_24_payload      ), //i
    .keyStatus_25_valid    (clk50Area_hid_keyStatus_25_valid        ), //i
    .keyStatus_25_payload  (clk50Area_hid_keyStatus_25_payload      ), //i
    .keyStatus_26_valid    (clk50Area_hid_keyStatus_26_valid        ), //i
    .keyStatus_26_payload  (clk50Area_hid_keyStatus_26_payload      ), //i
    .keyStatus_27_valid    (clk50Area_hid_keyStatus_27_valid        ), //i
    .keyStatus_27_payload  (clk50Area_hid_keyStatus_27_payload      ), //i
    .keyStatus_28_valid    (clk50Area_hid_keyStatus_28_valid        ), //i
    .keyStatus_28_payload  (clk50Area_hid_keyStatus_28_payload      ), //i
    .keyStatus_29_valid    (clk50Area_hid_keyStatus_29_valid        ), //i
    .keyStatus_29_payload  (clk50Area_hid_keyStatus_29_payload      ), //i
    .keyStatus_30_valid    (clk50Area_hid_keyStatus_30_valid        ), //i
    .keyStatus_30_payload  (clk50Area_hid_keyStatus_30_payload      ), //i
    .keyStatus_31_valid    (clk50Area_hid_keyStatus_31_valid        ), //i
    .keyStatus_31_payload  (clk50Area_hid_keyStatus_31_payload      ), //i
    .keyStatus_32_valid    (clk50Area_hid_keyStatus_32_valid        ), //i
    .keyStatus_32_payload  (clk50Area_hid_keyStatus_32_payload      ), //i
    .keyStatus_33_valid    (clk50Area_hid_keyStatus_33_valid        ), //i
    .keyStatus_33_payload  (clk50Area_hid_keyStatus_33_payload      ), //i
    .keyStatus_34_valid    (clk50Area_hid_keyStatus_34_valid        ), //i
    .keyStatus_34_payload  (clk50Area_hid_keyStatus_34_payload      ), //i
    .keyStatus_35_valid    (clk50Area_hid_keyStatus_35_valid        ), //i
    .keyStatus_35_payload  (clk50Area_hid_keyStatus_35_payload      ), //i
    .keyStatus_36_valid    (clk50Area_hid_keyStatus_36_valid        ), //i
    .keyStatus_36_payload  (clk50Area_hid_keyStatus_36_payload      ), //i
    .keyStatus_37_valid    (clk50Area_hid_keyStatus_37_valid        ), //i
    .keyStatus_37_payload  (clk50Area_hid_keyStatus_37_payload      ), //i
    .keyStatus_38_valid    (clk50Area_hid_keyStatus_38_valid        ), //i
    .keyStatus_38_payload  (clk50Area_hid_keyStatus_38_payload      ), //i
    .keyStatus_39_valid    (clk50Area_hid_keyStatus_39_valid        ), //i
    .keyStatus_39_payload  (clk50Area_hid_keyStatus_39_payload      ), //i
    .keyStatus_40_valid    (clk50Area_hid_keyStatus_40_valid        ), //i
    .keyStatus_40_payload  (clk50Area_hid_keyStatus_40_payload      ), //i
    .keyStatus_41_valid    (clk50Area_hid_keyStatus_41_valid        ), //i
    .keyStatus_41_payload  (clk50Area_hid_keyStatus_41_payload      ), //i
    .keyStatus_42_valid    (clk50Area_hid_keyStatus_42_valid        ), //i
    .keyStatus_42_payload  (clk50Area_hid_keyStatus_42_payload      ), //i
    .keyStatus_43_valid    (clk50Area_hid_keyStatus_43_valid        ), //i
    .keyStatus_43_payload  (clk50Area_hid_keyStatus_43_payload      ), //i
    .keyStatus_44_valid    (clk50Area_hid_keyStatus_44_valid        ), //i
    .keyStatus_44_payload  (clk50Area_hid_keyStatus_44_payload      ), //i
    .keyStatus_45_valid    (clk50Area_hid_keyStatus_45_valid        ), //i
    .keyStatus_45_payload  (clk50Area_hid_keyStatus_45_payload      ), //i
    .keyStatus_46_valid    (clk50Area_hid_keyStatus_46_valid        ), //i
    .keyStatus_46_payload  (clk50Area_hid_keyStatus_46_payload      ), //i
    .keyStatus_47_valid    (clk50Area_hid_keyStatus_47_valid        ), //i
    .keyStatus_47_payload  (clk50Area_hid_keyStatus_47_payload      ), //i
    .keyStatus_48_valid    (clk50Area_hid_keyStatus_48_valid        ), //i
    .keyStatus_48_payload  (clk50Area_hid_keyStatus_48_payload      ), //i
    .keyStatus_49_valid    (clk50Area_hid_keyStatus_49_valid        ), //i
    .keyStatus_49_payload  (clk50Area_hid_keyStatus_49_payload      ), //i
    .keyStatus_50_valid    (clk50Area_hid_keyStatus_50_valid        ), //i
    .keyStatus_50_payload  (clk50Area_hid_keyStatus_50_payload      ), //i
    .keyStatus_51_valid    (clk50Area_hid_keyStatus_51_valid        ), //i
    .keyStatus_51_payload  (clk50Area_hid_keyStatus_51_payload      ), //i
    .keyStatus_52_valid    (clk50Area_hid_keyStatus_52_valid        ), //i
    .keyStatus_52_payload  (clk50Area_hid_keyStatus_52_payload      ), //i
    .keyStatus_53_valid    (clk50Area_hid_keyStatus_53_valid        ), //i
    .keyStatus_53_payload  (clk50Area_hid_keyStatus_53_payload      ), //i
    .keyStatus_54_valid    (clk50Area_hid_keyStatus_54_valid        ), //i
    .keyStatus_54_payload  (clk50Area_hid_keyStatus_54_payload      ), //i
    .keyStatus_55_valid    (clk50Area_hid_keyStatus_55_valid        ), //i
    .keyStatus_55_payload  (clk50Area_hid_keyStatus_55_payload      ), //i
    .keyStatus_56_valid    (clk50Area_hid_keyStatus_56_valid        ), //i
    .keyStatus_56_payload  (clk50Area_hid_keyStatus_56_payload      ), //i
    .keyStatus_57_valid    (clk50Area_hid_keyStatus_57_valid        ), //i
    .keyStatus_57_payload  (clk50Area_hid_keyStatus_57_payload      ), //i
    .keyStatus_58_valid    (clk50Area_hid_keyStatus_58_valid        ), //i
    .keyStatus_58_payload  (clk50Area_hid_keyStatus_58_payload      ), //i
    .keyStatus_59_valid    (clk50Area_hid_keyStatus_59_valid        ), //i
    .keyStatus_59_payload  (clk50Area_hid_keyStatus_59_payload      ), //i
    .keyStatus_60_valid    (clk50Area_hid_keyStatus_60_valid        ), //i
    .keyStatus_60_payload  (clk50Area_hid_keyStatus_60_payload      ), //i
    .keyStatus_61_valid    (clk50Area_hid_keyStatus_61_valid        ), //i
    .keyStatus_61_payload  (clk50Area_hid_keyStatus_61_payload      ), //i
    .keyStatus_62_valid    (clk50Area_hid_keyStatus_62_valid        ), //i
    .keyStatus_62_payload  (clk50Area_hid_keyStatus_62_payload      ), //i
    .keyStatus_63_valid    (clk50Area_hid_keyStatus_63_valid        ), //i
    .keyStatus_63_payload  (clk50Area_hid_keyStatus_63_payload      ), //i
    .keyStatus_64_valid    (clk50Area_hid_keyStatus_64_valid        ), //i
    .keyStatus_64_payload  (clk50Area_hid_keyStatus_64_payload      ), //i
    .keyStatus_65_valid    (clk50Area_hid_keyStatus_65_valid        ), //i
    .keyStatus_65_payload  (clk50Area_hid_keyStatus_65_payload      ), //i
    .keyStatus_66_valid    (clk50Area_hid_keyStatus_66_valid        ), //i
    .keyStatus_66_payload  (clk50Area_hid_keyStatus_66_payload      ), //i
    .keyStatus_67_valid    (clk50Area_hid_keyStatus_67_valid        ), //i
    .keyStatus_67_payload  (clk50Area_hid_keyStatus_67_payload      ), //i
    .keyStatus_68_valid    (clk50Area_hid_keyStatus_68_valid        ), //i
    .keyStatus_68_payload  (clk50Area_hid_keyStatus_68_payload      ), //i
    .keyStatus_69_valid    (clk50Area_hid_keyStatus_69_valid        ), //i
    .keyStatus_69_payload  (clk50Area_hid_keyStatus_69_payload      ), //i
    .keyStatus_70_valid    (clk50Area_hid_keyStatus_70_valid        ), //i
    .keyStatus_70_payload  (clk50Area_hid_keyStatus_70_payload      ), //i
    .keyStatus_71_valid    (clk50Area_hid_keyStatus_71_valid        ), //i
    .keyStatus_71_payload  (clk50Area_hid_keyStatus_71_payload      ), //i
    .keyStatus_72_valid    (clk50Area_hid_keyStatus_72_valid        ), //i
    .keyStatus_72_payload  (clk50Area_hid_keyStatus_72_payload      ), //i
    .keyStatus_73_valid    (clk50Area_hid_keyStatus_73_valid        ), //i
    .keyStatus_73_payload  (clk50Area_hid_keyStatus_73_payload      ), //i
    .keyStatus_74_valid    (clk50Area_keyMatrix_keyStatus_74_valid  ), //i
    .keyStatus_74_payload  (clk50Area_keyMatrix_keyStatus_74_payload), //i
    .keyStatus_75_valid    (clk50Area_hid_keyStatus_75_valid        ), //i
    .keyStatus_75_payload  (clk50Area_hid_keyStatus_75_payload      ), //i
    .keyStatus_76_valid    (clk50Area_hid_keyStatus_76_valid        ), //i
    .keyStatus_76_payload  (clk50Area_hid_keyStatus_76_payload      ), //i
    .keyStatus_77_valid    (clk50Area_hid_keyStatus_77_valid        ), //i
    .keyStatus_77_payload  (clk50Area_hid_keyStatus_77_payload      ), //i
    .keyStatus_78_valid    (clk50Area_hid_keyStatus_78_valid        ), //i
    .keyStatus_78_payload  (clk50Area_hid_keyStatus_78_payload      ), //i
    .keyStatus_79_valid    (clk50Area_hid_keyStatus_79_valid        ), //i
    .keyStatus_79_payload  (clk50Area_hid_keyStatus_79_payload      ), //i
    .keyStatus_80_valid    (clk50Area_hid_keyStatus_80_valid        ), //i
    .keyStatus_80_payload  (clk50Area_hid_keyStatus_80_payload      ), //i
    .keyStatus_81_valid    (clk50Area_hid_keyStatus_81_valid        ), //i
    .keyStatus_81_payload  (clk50Area_hid_keyStatus_81_payload      ), //i
    .keyStatus_82_valid    (clk50Area_hid_keyStatus_82_valid        ), //i
    .keyStatus_82_payload  (clk50Area_hid_keyStatus_82_payload      ), //i
    .keyStatus_83_valid    (clk50Area_hid_keyStatus_83_valid        ), //i
    .keyStatus_83_payload  (clk50Area_hid_keyStatus_83_payload      ), //i
    .keyStatus_84_valid    (clk50Area_hid_keyStatus_84_valid        ), //i
    .keyStatus_84_payload  (clk50Area_hid_keyStatus_84_payload      ), //i
    .keyStatus_85_valid    (clk50Area_keyMatrix_keyStatus_85_valid  ), //i
    .keyStatus_85_payload  (clk50Area_keyMatrix_keyStatus_85_payload), //i
    .keyStatus_86_valid    (clk50Area_hid_keyStatus_86_valid        ), //i
    .keyStatus_86_payload  (clk50Area_hid_keyStatus_86_payload      ), //i
    .keyStatus_87_valid    (clk50Area_hid_keyStatus_87_valid        ), //i
    .keyStatus_87_payload  (clk50Area_hid_keyStatus_87_payload      ), //i
    .keyStatus_88_valid    (clk50Area_hid_keyStatus_88_valid        ), //i
    .keyStatus_88_payload  (clk50Area_hid_keyStatus_88_payload      ), //i
    .keyStatus_89_valid    (clk50Area_hid_keyStatus_89_valid        ), //i
    .keyStatus_89_payload  (clk50Area_hid_keyStatus_89_payload      ), //i
    .keyStatus_90_valid    (clk50Area_keyMatrix_keyStatus_90_valid  ), //i
    .keyStatus_90_payload  (clk50Area_keyMatrix_keyStatus_90_payload), //i
    .keyStatus_91_valid    (clk50Area_keyMatrix_keyStatus_91_valid  ), //i
    .keyStatus_91_payload  (clk50Area_keyMatrix_keyStatus_91_payload), //i
    .keyStatus_92_valid    (clk50Area_keyMatrix_keyStatus_92_valid  ), //i
    .keyStatus_92_payload  (clk50Area_keyMatrix_keyStatus_92_payload), //i
    .keyStatus_93_valid    (clk50Area_hid_keyStatus_93_valid        ), //i
    .keyStatus_93_payload  (clk50Area_hid_keyStatus_93_payload      ), //i
    .keyStatus_94_valid    (clk50Area_keyMatrix_keyStatus_94_valid  ), //i
    .keyStatus_94_payload  (clk50Area_keyMatrix_keyStatus_94_payload), //i
    .keyStatus_95_valid    (clk50Area_hid_keyStatus_95_valid        ), //i
    .keyStatus_95_payload  (clk50Area_hid_keyStatus_95_payload      ), //i
    .keyStatus_96_valid    (clk50Area_keyMatrix_keyStatus_96_valid  ), //i
    .keyStatus_96_payload  (clk50Area_keyMatrix_keyStatus_96_payload), //i
    .keyStatus_97_valid    (clk50Area_hid_keyStatus_97_valid        ), //i
    .keyStatus_97_payload  (clk50Area_hid_keyStatus_97_payload      ), //i
    .keyStatus_98_valid    (clk50Area_hid_keyStatus_98_valid        ), //i
    .keyStatus_98_payload  (clk50Area_hid_keyStatus_98_payload      ), //i
    .keyStatus_99_valid    (clk50Area_hid_keyStatus_99_valid        ), //i
    .keyStatus_99_payload  (clk50Area_hid_keyStatus_99_payload      ), //i
    .keyStatus_100_valid   (clk50Area_hid_keyStatus_100_valid       ), //i
    .keyStatus_100_payload (clk50Area_hid_keyStatus_100_payload     ), //i
    .keyStatus_101_valid   (clk50Area_hid_keyStatus_101_valid       ), //i
    .keyStatus_101_payload (clk50Area_hid_keyStatus_101_payload     ), //i
    .keyStatus_102_valid   (clk50Area_hid_keyStatus_102_valid       ), //i
    .keyStatus_102_payload (clk50Area_hid_keyStatus_102_payload     ), //i
    .CLK_50                (CLK_50                                  ), //i
    ._zz_LED_R6            (_zz_LED_R6                              )  //i
  );
  assign rstCtrl_io_externalReset = (! KEY_Fn);
  always @(*) begin
    _zz_LED_R6 = 1'b0;
    _zz_LED_R6 = bufferCC_3_io_dataOut;
  end

  assign _zz_1 = (rstCtrl_io_globalReset || (! pll100_locked));
  assign core_reset_reset_n = (! _zz_LED_R6);
  assign LED_A = core_io_row;
  assign LED_K = core_io_col;
  assign flash_dclk = core_flash_dclk;
  assign flash_sce = core_flash_sce;
  assign flash_sdo = core_flash_sdo;
  assign LED_R6 = _zz_LED_R6;
  assign ROW = clk50Area_keyMatrix_ROW;
  assign TXD = clk50Area_hid_TXD;
  always @(posedge CLK_50) begin
    if(clk50Area_keyMatrix_scanIdx_valid) begin
      toplevel_clk50Area_keyMatrix_scanIdx_payload_regNextWhen <= clk50Area_keyMatrix_scanIdx_payload;
    end
  end

  always @(posedge CLK_50 or posedge _zz_LED_R6) begin
    if(_zz_LED_R6) begin
      _zz_io_write_valid <= 1'b0;
    end else begin
      if(clk50Area_keyMatrix_scanIdx_valid) begin
        _zz_io_write_valid <= 1'b1;
      end else begin
        if(uartCtrl_2_io_write_ready) begin
          _zz_io_write_valid <= 1'b0;
        end
      end
    end
  end


endmodule

module HID (
  output              TXD,
  input               scanIdx_valid,
  input      [7:0]    scanIdx_payload,
  input               keyStatus_0_valid,
  input               keyStatus_0_payload,
  input               keyStatus_1_valid,
  input               keyStatus_1_payload,
  input               keyStatus_2_valid,
  input               keyStatus_2_payload,
  input               keyStatus_3_valid,
  input               keyStatus_3_payload,
  input               keyStatus_4_valid,
  input               keyStatus_4_payload,
  input               keyStatus_5_valid,
  input               keyStatus_5_payload,
  input               keyStatus_6_valid,
  input               keyStatus_6_payload,
  input               keyStatus_7_valid,
  input               keyStatus_7_payload,
  input               keyStatus_8_valid,
  input               keyStatus_8_payload,
  input               keyStatus_9_valid,
  input               keyStatus_9_payload,
  input               keyStatus_10_valid,
  input               keyStatus_10_payload,
  input               keyStatus_11_valid,
  input               keyStatus_11_payload,
  input               keyStatus_12_valid,
  input               keyStatus_12_payload,
  input               keyStatus_13_valid,
  input               keyStatus_13_payload,
  input               keyStatus_14_valid,
  input               keyStatus_14_payload,
  input               keyStatus_15_valid,
  input               keyStatus_15_payload,
  input               keyStatus_16_valid,
  input               keyStatus_16_payload,
  input               keyStatus_17_valid,
  input               keyStatus_17_payload,
  input               keyStatus_18_valid,
  input               keyStatus_18_payload,
  input               keyStatus_19_valid,
  input               keyStatus_19_payload,
  input               keyStatus_20_valid,
  input               keyStatus_20_payload,
  input               keyStatus_21_valid,
  input               keyStatus_21_payload,
  input               keyStatus_22_valid,
  input               keyStatus_22_payload,
  input               keyStatus_23_valid,
  input               keyStatus_23_payload,
  input               keyStatus_24_valid,
  input               keyStatus_24_payload,
  input               keyStatus_25_valid,
  input               keyStatus_25_payload,
  input               keyStatus_26_valid,
  input               keyStatus_26_payload,
  input               keyStatus_27_valid,
  input               keyStatus_27_payload,
  input               keyStatus_28_valid,
  input               keyStatus_28_payload,
  input               keyStatus_29_valid,
  input               keyStatus_29_payload,
  input               keyStatus_30_valid,
  input               keyStatus_30_payload,
  input               keyStatus_31_valid,
  input               keyStatus_31_payload,
  input               keyStatus_32_valid,
  input               keyStatus_32_payload,
  input               keyStatus_33_valid,
  input               keyStatus_33_payload,
  input               keyStatus_34_valid,
  input               keyStatus_34_payload,
  input               keyStatus_35_valid,
  input               keyStatus_35_payload,
  input               keyStatus_36_valid,
  input               keyStatus_36_payload,
  input               keyStatus_37_valid,
  input               keyStatus_37_payload,
  input               keyStatus_38_valid,
  input               keyStatus_38_payload,
  input               keyStatus_39_valid,
  input               keyStatus_39_payload,
  input               keyStatus_40_valid,
  input               keyStatus_40_payload,
  input               keyStatus_41_valid,
  input               keyStatus_41_payload,
  input               keyStatus_42_valid,
  input               keyStatus_42_payload,
  input               keyStatus_43_valid,
  input               keyStatus_43_payload,
  input               keyStatus_44_valid,
  input               keyStatus_44_payload,
  input               keyStatus_45_valid,
  input               keyStatus_45_payload,
  input               keyStatus_46_valid,
  input               keyStatus_46_payload,
  input               keyStatus_47_valid,
  input               keyStatus_47_payload,
  input               keyStatus_48_valid,
  input               keyStatus_48_payload,
  input               keyStatus_49_valid,
  input               keyStatus_49_payload,
  input               keyStatus_50_valid,
  input               keyStatus_50_payload,
  input               keyStatus_51_valid,
  input               keyStatus_51_payload,
  input               keyStatus_52_valid,
  input               keyStatus_52_payload,
  input               keyStatus_53_valid,
  input               keyStatus_53_payload,
  input               keyStatus_54_valid,
  input               keyStatus_54_payload,
  input               keyStatus_55_valid,
  input               keyStatus_55_payload,
  input               keyStatus_56_valid,
  input               keyStatus_56_payload,
  input               keyStatus_57_valid,
  input               keyStatus_57_payload,
  input               keyStatus_58_valid,
  input               keyStatus_58_payload,
  input               keyStatus_59_valid,
  input               keyStatus_59_payload,
  input               keyStatus_60_valid,
  input               keyStatus_60_payload,
  input               keyStatus_61_valid,
  input               keyStatus_61_payload,
  input               keyStatus_62_valid,
  input               keyStatus_62_payload,
  input               keyStatus_63_valid,
  input               keyStatus_63_payload,
  input               keyStatus_64_valid,
  input               keyStatus_64_payload,
  input               keyStatus_65_valid,
  input               keyStatus_65_payload,
  input               keyStatus_66_valid,
  input               keyStatus_66_payload,
  input               keyStatus_67_valid,
  input               keyStatus_67_payload,
  input               keyStatus_68_valid,
  input               keyStatus_68_payload,
  input               keyStatus_69_valid,
  input               keyStatus_69_payload,
  input               keyStatus_70_valid,
  input               keyStatus_70_payload,
  input               keyStatus_71_valid,
  input               keyStatus_71_payload,
  input               keyStatus_72_valid,
  input               keyStatus_72_payload,
  input               keyStatus_73_valid,
  input               keyStatus_73_payload,
  input               keyStatus_74_valid,
  input               keyStatus_74_payload,
  input               keyStatus_75_valid,
  input               keyStatus_75_payload,
  input               keyStatus_76_valid,
  input               keyStatus_76_payload,
  input               keyStatus_77_valid,
  input               keyStatus_77_payload,
  input               keyStatus_78_valid,
  input               keyStatus_78_payload,
  input               keyStatus_79_valid,
  input               keyStatus_79_payload,
  input               keyStatus_80_valid,
  input               keyStatus_80_payload,
  input               keyStatus_81_valid,
  input               keyStatus_81_payload,
  input               keyStatus_82_valid,
  input               keyStatus_82_payload,
  input               keyStatus_83_valid,
  input               keyStatus_83_payload,
  input               keyStatus_84_valid,
  input               keyStatus_84_payload,
  input               keyStatus_85_valid,
  input               keyStatus_85_payload,
  input               keyStatus_86_valid,
  input               keyStatus_86_payload,
  input               keyStatus_87_valid,
  input               keyStatus_87_payload,
  input               keyStatus_88_valid,
  input               keyStatus_88_payload,
  input               keyStatus_89_valid,
  input               keyStatus_89_payload,
  input               keyStatus_90_valid,
  input               keyStatus_90_payload,
  input               keyStatus_91_valid,
  input               keyStatus_91_payload,
  input               keyStatus_92_valid,
  input               keyStatus_92_payload,
  input               keyStatus_93_valid,
  input               keyStatus_93_payload,
  input               keyStatus_94_valid,
  input               keyStatus_94_payload,
  input               keyStatus_95_valid,
  input               keyStatus_95_payload,
  input               keyStatus_96_valid,
  input               keyStatus_96_payload,
  input               keyStatus_97_valid,
  input               keyStatus_97_payload,
  input               keyStatus_98_valid,
  input               keyStatus_98_payload,
  input               keyStatus_99_valid,
  input               keyStatus_99_payload,
  input               keyStatus_100_valid,
  input               keyStatus_100_payload,
  input               keyStatus_101_valid,
  input               keyStatus_101_payload,
  input               keyStatus_102_valid,
  input               keyStatus_102_payload,
  input               CLK_50,
  input               _zz_LED_R6
);
  localparam UartParityType_NONE = 2'd0;
  localparam UartParityType_EVEN = 2'd1;
  localparam UartParityType_ODD = 2'd2;
  localparam UartStopType_ONE = 1'd0;
  localparam UartStopType_TWO = 1'd1;
  localparam machine_enumDef_BOOT = 4'd0;
  localparam machine_enumDef_idle = 4'd1;
  localparam machine_enumDef_k6 = 4'd2;
  localparam machine_enumDef_k5 = 4'd3;
  localparam machine_enumDef_k4 = 4'd4;
  localparam machine_enumDef_k3 = 4'd5;
  localparam machine_enumDef_k2 = 4'd6;
  localparam machine_enumDef_k1 = 4'd7;
  localparam machine_enumDef_reserved = 4'd8;
  localparam machine_enumDef_special = 4'd9;

  wire                uartCtrl_2_io_write_valid;
  reg        [7:0]    uartCtrl_2_io_write_payload;
  wire                uartCtrl_2_io_read_ready;
  reg        [7:0]    _zz_hidKeyTable_port0;
  wire                uartCtrl_2_io_write_ready;
  wire                uartCtrl_2_io_read_valid;
  wire       [7:0]    uartCtrl_2_io_read_payload;
  wire                uartCtrl_2_io_uart_txd;
  wire                uartCtrl_2_io_readError;
  wire                uartCtrl_2_io_readBreak;
  wire                _zz_hidKeyTable_port;
  wire                _zz_io_write_payload;
  reg        [6:0]    idxLatch;
  reg                 staLatch;
  wire                machine_wantExit;
  reg                 machine_wantStart;
  wire                machine_wantKill;
  reg        [3:0]    machine_stateReg;
  reg        [3:0]    machine_stateNext;
  `ifndef SYNTHESIS
  reg [63:0] machine_stateReg_string;
  reg [63:0] machine_stateNext_string;
  `endif

  (* ram_init_file = "VerilogHDL/hid.mif" *) reg [7:0] hidKeyTable [0:127];

  assign _zz_io_write_payload = 1'b1;
  always @(posedge CLK_50) begin
    if(_zz_io_write_payload) begin
      _zz_hidKeyTable_port0 <= hidKeyTable[idxLatch];
    end
  end

  UartCtrl_1 uartCtrl_2 (
    .io_config_frame_dataLength (3'b111                          ), //i
    .io_config_frame_stop       (UartStopType_ONE                ), //i
    .io_config_frame_parity     (UartParityType_NONE             ), //i
    .io_config_clockDivider     (20'h0028a                       ), //i
    .io_write_valid             (uartCtrl_2_io_write_valid       ), //i
    .io_write_ready             (uartCtrl_2_io_write_ready       ), //o
    .io_write_payload           (uartCtrl_2_io_write_payload[7:0]), //i
    .io_read_valid              (uartCtrl_2_io_read_valid        ), //o
    .io_read_ready              (uartCtrl_2_io_read_ready        ), //i
    .io_read_payload            (uartCtrl_2_io_read_payload[7:0] ), //o
    .io_uart_txd                (uartCtrl_2_io_uart_txd          ), //o
    .io_uart_rxd                (1'b1                            ), //i
    .io_readError               (uartCtrl_2_io_readError         ), //o
    .io_writeBreak              (1'b0                            ), //i
    .io_readBreak               (uartCtrl_2_io_readBreak         ), //o
    .CLK_50                     (CLK_50                          ), //i
    ._zz_LED_R6                 (_zz_LED_R6                      )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(machine_stateReg)
      machine_enumDef_BOOT : machine_stateReg_string = "BOOT    ";
      machine_enumDef_idle : machine_stateReg_string = "idle    ";
      machine_enumDef_k6 : machine_stateReg_string = "k6      ";
      machine_enumDef_k5 : machine_stateReg_string = "k5      ";
      machine_enumDef_k4 : machine_stateReg_string = "k4      ";
      machine_enumDef_k3 : machine_stateReg_string = "k3      ";
      machine_enumDef_k2 : machine_stateReg_string = "k2      ";
      machine_enumDef_k1 : machine_stateReg_string = "k1      ";
      machine_enumDef_reserved : machine_stateReg_string = "reserved";
      machine_enumDef_special : machine_stateReg_string = "special ";
      default : machine_stateReg_string = "????????";
    endcase
  end
  always @(*) begin
    case(machine_stateNext)
      machine_enumDef_BOOT : machine_stateNext_string = "BOOT    ";
      machine_enumDef_idle : machine_stateNext_string = "idle    ";
      machine_enumDef_k6 : machine_stateNext_string = "k6      ";
      machine_enumDef_k5 : machine_stateNext_string = "k5      ";
      machine_enumDef_k4 : machine_stateNext_string = "k4      ";
      machine_enumDef_k3 : machine_stateNext_string = "k3      ";
      machine_enumDef_k2 : machine_stateNext_string = "k2      ";
      machine_enumDef_k1 : machine_stateNext_string = "k1      ";
      machine_enumDef_reserved : machine_stateNext_string = "reserved";
      machine_enumDef_special : machine_stateNext_string = "special ";
      default : machine_stateNext_string = "????????";
    endcase
  end
  `endif

  always @(*) begin
    uartCtrl_2_io_write_payload = 8'h0;
    case(machine_stateReg)
      machine_enumDef_idle : begin
      end
      machine_enumDef_k6 : begin
      end
      machine_enumDef_k5 : begin
      end
      machine_enumDef_k4 : begin
      end
      machine_enumDef_k3 : begin
      end
      machine_enumDef_k2 : begin
      end
      machine_enumDef_k1 : begin
        if(staLatch) begin
          uartCtrl_2_io_write_payload = _zz_hidKeyTable_port0;
        end
      end
      machine_enumDef_reserved : begin
      end
      machine_enumDef_special : begin
        uartCtrl_2_io_write_payload = {1'b0,{keyStatus_94_payload,{keyStatus_85_payload,{keyStatus_96_payload,{keyStatus_91_payload,{keyStatus_92_payload,{keyStatus_74_payload,keyStatus_90_payload}}}}}}};
      end
      default : begin
      end
    endcase
  end

  assign TXD = uartCtrl_2_io_uart_txd;
  assign machine_wantExit = 1'b0;
  always @(*) begin
    machine_wantStart = 1'b0;
    case(machine_stateReg)
      machine_enumDef_idle : begin
      end
      machine_enumDef_k6 : begin
      end
      machine_enumDef_k5 : begin
      end
      machine_enumDef_k4 : begin
      end
      machine_enumDef_k3 : begin
      end
      machine_enumDef_k2 : begin
      end
      machine_enumDef_k1 : begin
      end
      machine_enumDef_reserved : begin
      end
      machine_enumDef_special : begin
      end
      default : begin
        machine_wantStart = 1'b1;
      end
    endcase
  end

  assign machine_wantKill = 1'b0;
  assign uartCtrl_2_io_write_valid = (! (machine_stateReg == machine_enumDef_idle));
  always @(*) begin
    machine_stateNext = machine_stateReg;
    case(machine_stateReg)
      machine_enumDef_idle : begin
        if(scanIdx_valid) begin
          machine_stateNext = machine_enumDef_special;
        end
      end
      machine_enumDef_k6 : begin
        if(uartCtrl_2_io_write_ready) begin
          machine_stateNext = machine_enumDef_idle;
        end
      end
      machine_enumDef_k5 : begin
        if(uartCtrl_2_io_write_ready) begin
          machine_stateNext = machine_enumDef_k6;
        end
      end
      machine_enumDef_k4 : begin
        if(uartCtrl_2_io_write_ready) begin
          machine_stateNext = machine_enumDef_k5;
        end
      end
      machine_enumDef_k3 : begin
        if(uartCtrl_2_io_write_ready) begin
          machine_stateNext = machine_enumDef_k4;
        end
      end
      machine_enumDef_k2 : begin
        if(uartCtrl_2_io_write_ready) begin
          machine_stateNext = machine_enumDef_k3;
        end
      end
      machine_enumDef_k1 : begin
        if(uartCtrl_2_io_write_ready) begin
          machine_stateNext = machine_enumDef_k2;
        end
      end
      machine_enumDef_reserved : begin
        if(uartCtrl_2_io_write_ready) begin
          machine_stateNext = machine_enumDef_k1;
        end
      end
      machine_enumDef_special : begin
        if(uartCtrl_2_io_write_ready) begin
          machine_stateNext = machine_enumDef_reserved;
        end
      end
      default : begin
      end
    endcase
    if(machine_wantStart) begin
      machine_stateNext = machine_enumDef_idle;
    end
    if(machine_wantKill) begin
      machine_stateNext = machine_enumDef_BOOT;
    end
  end

  always @(posedge CLK_50 or posedge _zz_LED_R6) begin
    if(_zz_LED_R6) begin
      idxLatch <= 7'h0;
      staLatch <= 1'b0;
      machine_stateReg <= machine_enumDef_BOOT;
    end else begin
      if(scanIdx_valid) begin
        idxLatch <= scanIdx_payload[6 : 0];
      end
      if(scanIdx_valid) begin
        staLatch <= scanIdx_payload[7];
      end
      machine_stateReg <= machine_stateNext;
    end
  end


endmodule

//UartCtrl_1 replaced by UartCtrl_1

module KeyMatrix (
  input               enabled,
  input      [20:0]   COL,
  output     [5:0]    ROW,
  output              scanIdx_valid,
  output     [7:0]    scanIdx_payload,
  output              keyStatus_0_valid,
  output              keyStatus_0_payload,
  output              keyStatus_1_valid,
  output              keyStatus_1_payload,
  output              keyStatus_2_valid,
  output              keyStatus_2_payload,
  output              keyStatus_3_valid,
  output              keyStatus_3_payload,
  output              keyStatus_4_valid,
  output              keyStatus_4_payload,
  output              keyStatus_5_valid,
  output              keyStatus_5_payload,
  output              keyStatus_6_valid,
  output              keyStatus_6_payload,
  output              keyStatus_7_valid,
  output              keyStatus_7_payload,
  output              keyStatus_8_valid,
  output              keyStatus_8_payload,
  output              keyStatus_9_valid,
  output              keyStatus_9_payload,
  output              keyStatus_10_valid,
  output              keyStatus_10_payload,
  output              keyStatus_11_valid,
  output              keyStatus_11_payload,
  output              keyStatus_12_valid,
  output              keyStatus_12_payload,
  output              keyStatus_13_valid,
  output              keyStatus_13_payload,
  output              keyStatus_14_valid,
  output              keyStatus_14_payload,
  output              keyStatus_15_valid,
  output              keyStatus_15_payload,
  output              keyStatus_16_valid,
  output              keyStatus_16_payload,
  output              keyStatus_17_valid,
  output              keyStatus_17_payload,
  output              keyStatus_18_valid,
  output              keyStatus_18_payload,
  output              keyStatus_19_valid,
  output              keyStatus_19_payload,
  output              keyStatus_20_valid,
  output              keyStatus_20_payload,
  output              keyStatus_21_valid,
  output              keyStatus_21_payload,
  output              keyStatus_22_valid,
  output              keyStatus_22_payload,
  output              keyStatus_23_valid,
  output              keyStatus_23_payload,
  output              keyStatus_24_valid,
  output              keyStatus_24_payload,
  output              keyStatus_25_valid,
  output              keyStatus_25_payload,
  output              keyStatus_26_valid,
  output              keyStatus_26_payload,
  output              keyStatus_27_valid,
  output              keyStatus_27_payload,
  output              keyStatus_28_valid,
  output              keyStatus_28_payload,
  output              keyStatus_29_valid,
  output              keyStatus_29_payload,
  output              keyStatus_30_valid,
  output              keyStatus_30_payload,
  output              keyStatus_31_valid,
  output              keyStatus_31_payload,
  output              keyStatus_32_valid,
  output              keyStatus_32_payload,
  output              keyStatus_33_valid,
  output              keyStatus_33_payload,
  output              keyStatus_34_valid,
  output              keyStatus_34_payload,
  output              keyStatus_35_valid,
  output              keyStatus_35_payload,
  output              keyStatus_36_valid,
  output              keyStatus_36_payload,
  output              keyStatus_37_valid,
  output              keyStatus_37_payload,
  output              keyStatus_38_valid,
  output              keyStatus_38_payload,
  output              keyStatus_39_valid,
  output              keyStatus_39_payload,
  output              keyStatus_40_valid,
  output              keyStatus_40_payload,
  output              keyStatus_41_valid,
  output              keyStatus_41_payload,
  output              keyStatus_42_valid,
  output              keyStatus_42_payload,
  output              keyStatus_43_valid,
  output              keyStatus_43_payload,
  output              keyStatus_44_valid,
  output              keyStatus_44_payload,
  output              keyStatus_45_valid,
  output              keyStatus_45_payload,
  output              keyStatus_46_valid,
  output              keyStatus_46_payload,
  output              keyStatus_47_valid,
  output              keyStatus_47_payload,
  output              keyStatus_48_valid,
  output              keyStatus_48_payload,
  output              keyStatus_49_valid,
  output              keyStatus_49_payload,
  output              keyStatus_50_valid,
  output              keyStatus_50_payload,
  output              keyStatus_51_valid,
  output              keyStatus_51_payload,
  output              keyStatus_52_valid,
  output              keyStatus_52_payload,
  output              keyStatus_53_valid,
  output              keyStatus_53_payload,
  output              keyStatus_54_valid,
  output              keyStatus_54_payload,
  output              keyStatus_55_valid,
  output              keyStatus_55_payload,
  output              keyStatus_56_valid,
  output              keyStatus_56_payload,
  output              keyStatus_57_valid,
  output              keyStatus_57_payload,
  output              keyStatus_58_valid,
  output              keyStatus_58_payload,
  output              keyStatus_59_valid,
  output              keyStatus_59_payload,
  output              keyStatus_60_valid,
  output              keyStatus_60_payload,
  output              keyStatus_61_valid,
  output              keyStatus_61_payload,
  output              keyStatus_62_valid,
  output              keyStatus_62_payload,
  output              keyStatus_63_valid,
  output              keyStatus_63_payload,
  output              keyStatus_64_valid,
  output              keyStatus_64_payload,
  output              keyStatus_65_valid,
  output              keyStatus_65_payload,
  output              keyStatus_66_valid,
  output              keyStatus_66_payload,
  output              keyStatus_67_valid,
  output              keyStatus_67_payload,
  output              keyStatus_68_valid,
  output              keyStatus_68_payload,
  output              keyStatus_69_valid,
  output              keyStatus_69_payload,
  output              keyStatus_70_valid,
  output              keyStatus_70_payload,
  output              keyStatus_71_valid,
  output              keyStatus_71_payload,
  output              keyStatus_72_valid,
  output              keyStatus_72_payload,
  output              keyStatus_73_valid,
  output              keyStatus_73_payload,
  output              keyStatus_74_valid,
  output              keyStatus_74_payload,
  output              keyStatus_75_valid,
  output              keyStatus_75_payload,
  output              keyStatus_76_valid,
  output              keyStatus_76_payload,
  output              keyStatus_77_valid,
  output              keyStatus_77_payload,
  output              keyStatus_78_valid,
  output              keyStatus_78_payload,
  output              keyStatus_79_valid,
  output              keyStatus_79_payload,
  output              keyStatus_80_valid,
  output              keyStatus_80_payload,
  output              keyStatus_81_valid,
  output              keyStatus_81_payload,
  output              keyStatus_82_valid,
  output              keyStatus_82_payload,
  output              keyStatus_83_valid,
  output              keyStatus_83_payload,
  output              keyStatus_84_valid,
  output              keyStatus_84_payload,
  output              keyStatus_85_valid,
  output              keyStatus_85_payload,
  output              keyStatus_86_valid,
  output              keyStatus_86_payload,
  output              keyStatus_87_valid,
  output              keyStatus_87_payload,
  output              keyStatus_88_valid,
  output              keyStatus_88_payload,
  output              keyStatus_89_valid,
  output              keyStatus_89_payload,
  output              keyStatus_90_valid,
  output              keyStatus_90_payload,
  output              keyStatus_91_valid,
  output              keyStatus_91_payload,
  output              keyStatus_92_valid,
  output              keyStatus_92_payload,
  output              keyStatus_93_valid,
  output              keyStatus_93_payload,
  output              keyStatus_94_valid,
  output              keyStatus_94_payload,
  output              keyStatus_95_valid,
  output              keyStatus_95_payload,
  output              keyStatus_96_valid,
  output              keyStatus_96_payload,
  output              keyStatus_97_valid,
  output              keyStatus_97_payload,
  output              keyStatus_98_valid,
  output              keyStatus_98_payload,
  output              keyStatus_99_valid,
  output              keyStatus_99_payload,
  output              keyStatus_100_valid,
  output              keyStatus_100_payload,
  output              keyStatus_101_valid,
  output              keyStatus_101_payload,
  output              keyStatus_102_valid,
  output              keyStatus_102_payload,
  input               _zz_LED_R6,
  input               CLK_50
);

  wire       [5:0]    scanK_ROW;
  wire       [102:0]  scanK_key_down;
  wire                debounce_1_keyStatus_0_valid;
  wire                debounce_1_keyStatus_0_payload;
  wire                debounce_1_keyStatus_1_valid;
  wire                debounce_1_keyStatus_1_payload;
  wire                debounce_1_keyStatus_2_valid;
  wire                debounce_1_keyStatus_2_payload;
  wire                debounce_1_keyStatus_3_valid;
  wire                debounce_1_keyStatus_3_payload;
  wire                debounce_1_keyStatus_4_valid;
  wire                debounce_1_keyStatus_4_payload;
  wire                debounce_1_keyStatus_5_valid;
  wire                debounce_1_keyStatus_5_payload;
  wire                debounce_1_keyStatus_6_valid;
  wire                debounce_1_keyStatus_6_payload;
  wire                debounce_1_keyStatus_7_valid;
  wire                debounce_1_keyStatus_7_payload;
  wire                debounce_1_keyStatus_8_valid;
  wire                debounce_1_keyStatus_8_payload;
  wire                debounce_1_keyStatus_9_valid;
  wire                debounce_1_keyStatus_9_payload;
  wire                debounce_1_keyStatus_10_valid;
  wire                debounce_1_keyStatus_10_payload;
  wire                debounce_1_keyStatus_11_valid;
  wire                debounce_1_keyStatus_11_payload;
  wire                debounce_1_keyStatus_12_valid;
  wire                debounce_1_keyStatus_12_payload;
  wire                debounce_1_keyStatus_13_valid;
  wire                debounce_1_keyStatus_13_payload;
  wire                debounce_1_keyStatus_14_valid;
  wire                debounce_1_keyStatus_14_payload;
  wire                debounce_1_keyStatus_15_valid;
  wire                debounce_1_keyStatus_15_payload;
  wire                debounce_1_keyStatus_16_valid;
  wire                debounce_1_keyStatus_16_payload;
  wire                debounce_1_keyStatus_17_valid;
  wire                debounce_1_keyStatus_17_payload;
  wire                debounce_1_keyStatus_18_valid;
  wire                debounce_1_keyStatus_18_payload;
  wire                debounce_1_keyStatus_19_valid;
  wire                debounce_1_keyStatus_19_payload;
  wire                debounce_1_keyStatus_20_valid;
  wire                debounce_1_keyStatus_20_payload;
  wire                debounce_1_keyStatus_21_valid;
  wire                debounce_1_keyStatus_21_payload;
  wire                debounce_1_keyStatus_22_valid;
  wire                debounce_1_keyStatus_22_payload;
  wire                debounce_1_keyStatus_23_valid;
  wire                debounce_1_keyStatus_23_payload;
  wire                debounce_1_keyStatus_24_valid;
  wire                debounce_1_keyStatus_24_payload;
  wire                debounce_1_keyStatus_25_valid;
  wire                debounce_1_keyStatus_25_payload;
  wire                debounce_1_keyStatus_26_valid;
  wire                debounce_1_keyStatus_26_payload;
  wire                debounce_1_keyStatus_27_valid;
  wire                debounce_1_keyStatus_27_payload;
  wire                debounce_1_keyStatus_28_valid;
  wire                debounce_1_keyStatus_28_payload;
  wire                debounce_1_keyStatus_29_valid;
  wire                debounce_1_keyStatus_29_payload;
  wire                debounce_1_keyStatus_30_valid;
  wire                debounce_1_keyStatus_30_payload;
  wire                debounce_1_keyStatus_31_valid;
  wire                debounce_1_keyStatus_31_payload;
  wire                debounce_1_keyStatus_32_valid;
  wire                debounce_1_keyStatus_32_payload;
  wire                debounce_1_keyStatus_33_valid;
  wire                debounce_1_keyStatus_33_payload;
  wire                debounce_1_keyStatus_34_valid;
  wire                debounce_1_keyStatus_34_payload;
  wire                debounce_1_keyStatus_35_valid;
  wire                debounce_1_keyStatus_35_payload;
  wire                debounce_1_keyStatus_36_valid;
  wire                debounce_1_keyStatus_36_payload;
  wire                debounce_1_keyStatus_37_valid;
  wire                debounce_1_keyStatus_37_payload;
  wire                debounce_1_keyStatus_38_valid;
  wire                debounce_1_keyStatus_38_payload;
  wire                debounce_1_keyStatus_39_valid;
  wire                debounce_1_keyStatus_39_payload;
  wire                debounce_1_keyStatus_40_valid;
  wire                debounce_1_keyStatus_40_payload;
  wire                debounce_1_keyStatus_41_valid;
  wire                debounce_1_keyStatus_41_payload;
  wire                debounce_1_keyStatus_42_valid;
  wire                debounce_1_keyStatus_42_payload;
  wire                debounce_1_keyStatus_43_valid;
  wire                debounce_1_keyStatus_43_payload;
  wire                debounce_1_keyStatus_44_valid;
  wire                debounce_1_keyStatus_44_payload;
  wire                debounce_1_keyStatus_45_valid;
  wire                debounce_1_keyStatus_45_payload;
  wire                debounce_1_keyStatus_46_valid;
  wire                debounce_1_keyStatus_46_payload;
  wire                debounce_1_keyStatus_47_valid;
  wire                debounce_1_keyStatus_47_payload;
  wire                debounce_1_keyStatus_48_valid;
  wire                debounce_1_keyStatus_48_payload;
  wire                debounce_1_keyStatus_49_valid;
  wire                debounce_1_keyStatus_49_payload;
  wire                debounce_1_keyStatus_50_valid;
  wire                debounce_1_keyStatus_50_payload;
  wire                debounce_1_keyStatus_51_valid;
  wire                debounce_1_keyStatus_51_payload;
  wire                debounce_1_keyStatus_52_valid;
  wire                debounce_1_keyStatus_52_payload;
  wire                debounce_1_keyStatus_53_valid;
  wire                debounce_1_keyStatus_53_payload;
  wire                debounce_1_keyStatus_54_valid;
  wire                debounce_1_keyStatus_54_payload;
  wire                debounce_1_keyStatus_55_valid;
  wire                debounce_1_keyStatus_55_payload;
  wire                debounce_1_keyStatus_56_valid;
  wire                debounce_1_keyStatus_56_payload;
  wire                debounce_1_keyStatus_57_valid;
  wire                debounce_1_keyStatus_57_payload;
  wire                debounce_1_keyStatus_58_valid;
  wire                debounce_1_keyStatus_58_payload;
  wire                debounce_1_keyStatus_59_valid;
  wire                debounce_1_keyStatus_59_payload;
  wire                debounce_1_keyStatus_60_valid;
  wire                debounce_1_keyStatus_60_payload;
  wire                debounce_1_keyStatus_61_valid;
  wire                debounce_1_keyStatus_61_payload;
  wire                debounce_1_keyStatus_62_valid;
  wire                debounce_1_keyStatus_62_payload;
  wire                debounce_1_keyStatus_63_valid;
  wire                debounce_1_keyStatus_63_payload;
  wire                debounce_1_keyStatus_64_valid;
  wire                debounce_1_keyStatus_64_payload;
  wire                debounce_1_keyStatus_65_valid;
  wire                debounce_1_keyStatus_65_payload;
  wire                debounce_1_keyStatus_66_valid;
  wire                debounce_1_keyStatus_66_payload;
  wire                debounce_1_keyStatus_67_valid;
  wire                debounce_1_keyStatus_67_payload;
  wire                debounce_1_keyStatus_68_valid;
  wire                debounce_1_keyStatus_68_payload;
  wire                debounce_1_keyStatus_69_valid;
  wire                debounce_1_keyStatus_69_payload;
  wire                debounce_1_keyStatus_70_valid;
  wire                debounce_1_keyStatus_70_payload;
  wire                debounce_1_keyStatus_71_valid;
  wire                debounce_1_keyStatus_71_payload;
  wire                debounce_1_keyStatus_72_valid;
  wire                debounce_1_keyStatus_72_payload;
  wire                debounce_1_keyStatus_73_valid;
  wire                debounce_1_keyStatus_73_payload;
  wire                debounce_1_keyStatus_74_valid;
  wire                debounce_1_keyStatus_74_payload;
  wire                debounce_1_keyStatus_75_valid;
  wire                debounce_1_keyStatus_75_payload;
  wire                debounce_1_keyStatus_76_valid;
  wire                debounce_1_keyStatus_76_payload;
  wire                debounce_1_keyStatus_77_valid;
  wire                debounce_1_keyStatus_77_payload;
  wire                debounce_1_keyStatus_78_valid;
  wire                debounce_1_keyStatus_78_payload;
  wire                debounce_1_keyStatus_79_valid;
  wire                debounce_1_keyStatus_79_payload;
  wire                debounce_1_keyStatus_80_valid;
  wire                debounce_1_keyStatus_80_payload;
  wire                debounce_1_keyStatus_81_valid;
  wire                debounce_1_keyStatus_81_payload;
  wire                debounce_1_keyStatus_82_valid;
  wire                debounce_1_keyStatus_82_payload;
  wire                debounce_1_keyStatus_83_valid;
  wire                debounce_1_keyStatus_83_payload;
  wire                debounce_1_keyStatus_84_valid;
  wire                debounce_1_keyStatus_84_payload;
  wire                debounce_1_keyStatus_85_valid;
  wire                debounce_1_keyStatus_85_payload;
  wire                debounce_1_keyStatus_86_valid;
  wire                debounce_1_keyStatus_86_payload;
  wire                debounce_1_keyStatus_87_valid;
  wire                debounce_1_keyStatus_87_payload;
  wire                debounce_1_keyStatus_88_valid;
  wire                debounce_1_keyStatus_88_payload;
  wire                debounce_1_keyStatus_89_valid;
  wire                debounce_1_keyStatus_89_payload;
  wire                debounce_1_keyStatus_90_valid;
  wire                debounce_1_keyStatus_90_payload;
  wire                debounce_1_keyStatus_91_valid;
  wire                debounce_1_keyStatus_91_payload;
  wire                debounce_1_keyStatus_92_valid;
  wire                debounce_1_keyStatus_92_payload;
  wire                debounce_1_keyStatus_93_valid;
  wire                debounce_1_keyStatus_93_payload;
  wire                debounce_1_keyStatus_94_valid;
  wire                debounce_1_keyStatus_94_payload;
  wire                debounce_1_keyStatus_95_valid;
  wire                debounce_1_keyStatus_95_payload;
  wire                debounce_1_keyStatus_96_valid;
  wire                debounce_1_keyStatus_96_payload;
  wire                debounce_1_keyStatus_97_valid;
  wire                debounce_1_keyStatus_97_payload;
  wire                debounce_1_keyStatus_98_valid;
  wire                debounce_1_keyStatus_98_payload;
  wire                debounce_1_keyStatus_99_valid;
  wire                debounce_1_keyStatus_99_payload;
  wire                debounce_1_keyStatus_100_valid;
  wire                debounce_1_keyStatus_100_payload;
  wire                debounce_1_keyStatus_101_valid;
  wire                debounce_1_keyStatus_101_payload;
  wire                debounce_1_keyStatus_102_valid;
  wire                debounce_1_keyStatus_102_payload;
  wire       [12:0]   _zz_clkScan_counter_valueNext;
  wire       [0:0]    _zz_clkScan_counter_valueNext_1;
  wire       [6:0]    _zz__zz_scanIdx_valid_1;
  wire       [0:0]    _zz__zz_scanIdx_valid_1_1;
  reg                 _zz_scanIdx_valid_3;
  reg                 _zz_scanIdx_payload;
  reg                 clkScan_state;
  reg                 clkScan_stateRise;
  wire                clkScan_counter_willIncrement;
  reg                 clkScan_counter_willClear;
  reg        [12:0]   clkScan_counter_valueNext;
  reg        [12:0]   clkScan_counter_value;
  wire                clkScan_counter_willOverflowIfInc;
  wire                clkScan_counter_willOverflow;
  reg        [7:0]    _zz_when_ClockDomain_l369;
  wire                when_ClockDomain_l369;
  reg                 when_ClockDomain_l369_regNext;
  wire                _zz_scanIdx_valid;
  reg        [6:0]    _zz_scanIdx_valid_1;
  reg        [6:0]    _zz_scanIdx_valid_2;
  wire                _zz_1;
  wire                _zz_2;

  assign _zz_clkScan_counter_valueNext_1 = clkScan_counter_willIncrement;
  assign _zz_clkScan_counter_valueNext = {12'd0, _zz_clkScan_counter_valueNext_1};
  assign _zz__zz_scanIdx_valid_1_1 = _zz_scanIdx_valid;
  assign _zz__zz_scanIdx_valid_1 = {6'd0, _zz__zz_scanIdx_valid_1_1};
  scan_key scanK (
    .clock    (clkScan_state        ), //i
    .reset    (_zz_LED_R6           ), //i
    .enabled  (enabled              ), //i
    .COL      (COL[20:0]            ), //i
    .ROW      (scanK_ROW[5:0]       ), //o
    .key_down (scanK_key_down[102:0])  //o
  );
  Debounce debounce_1 (
    .key_down              (scanK_key_down[102:0]           ), //i
    .keyStatus_0_valid     (debounce_1_keyStatus_0_valid    ), //o
    .keyStatus_0_payload   (debounce_1_keyStatus_0_payload  ), //o
    .keyStatus_1_valid     (debounce_1_keyStatus_1_valid    ), //o
    .keyStatus_1_payload   (debounce_1_keyStatus_1_payload  ), //o
    .keyStatus_2_valid     (debounce_1_keyStatus_2_valid    ), //o
    .keyStatus_2_payload   (debounce_1_keyStatus_2_payload  ), //o
    .keyStatus_3_valid     (debounce_1_keyStatus_3_valid    ), //o
    .keyStatus_3_payload   (debounce_1_keyStatus_3_payload  ), //o
    .keyStatus_4_valid     (debounce_1_keyStatus_4_valid    ), //o
    .keyStatus_4_payload   (debounce_1_keyStatus_4_payload  ), //o
    .keyStatus_5_valid     (debounce_1_keyStatus_5_valid    ), //o
    .keyStatus_5_payload   (debounce_1_keyStatus_5_payload  ), //o
    .keyStatus_6_valid     (debounce_1_keyStatus_6_valid    ), //o
    .keyStatus_6_payload   (debounce_1_keyStatus_6_payload  ), //o
    .keyStatus_7_valid     (debounce_1_keyStatus_7_valid    ), //o
    .keyStatus_7_payload   (debounce_1_keyStatus_7_payload  ), //o
    .keyStatus_8_valid     (debounce_1_keyStatus_8_valid    ), //o
    .keyStatus_8_payload   (debounce_1_keyStatus_8_payload  ), //o
    .keyStatus_9_valid     (debounce_1_keyStatus_9_valid    ), //o
    .keyStatus_9_payload   (debounce_1_keyStatus_9_payload  ), //o
    .keyStatus_10_valid    (debounce_1_keyStatus_10_valid   ), //o
    .keyStatus_10_payload  (debounce_1_keyStatus_10_payload ), //o
    .keyStatus_11_valid    (debounce_1_keyStatus_11_valid   ), //o
    .keyStatus_11_payload  (debounce_1_keyStatus_11_payload ), //o
    .keyStatus_12_valid    (debounce_1_keyStatus_12_valid   ), //o
    .keyStatus_12_payload  (debounce_1_keyStatus_12_payload ), //o
    .keyStatus_13_valid    (debounce_1_keyStatus_13_valid   ), //o
    .keyStatus_13_payload  (debounce_1_keyStatus_13_payload ), //o
    .keyStatus_14_valid    (debounce_1_keyStatus_14_valid   ), //o
    .keyStatus_14_payload  (debounce_1_keyStatus_14_payload ), //o
    .keyStatus_15_valid    (debounce_1_keyStatus_15_valid   ), //o
    .keyStatus_15_payload  (debounce_1_keyStatus_15_payload ), //o
    .keyStatus_16_valid    (debounce_1_keyStatus_16_valid   ), //o
    .keyStatus_16_payload  (debounce_1_keyStatus_16_payload ), //o
    .keyStatus_17_valid    (debounce_1_keyStatus_17_valid   ), //o
    .keyStatus_17_payload  (debounce_1_keyStatus_17_payload ), //o
    .keyStatus_18_valid    (debounce_1_keyStatus_18_valid   ), //o
    .keyStatus_18_payload  (debounce_1_keyStatus_18_payload ), //o
    .keyStatus_19_valid    (debounce_1_keyStatus_19_valid   ), //o
    .keyStatus_19_payload  (debounce_1_keyStatus_19_payload ), //o
    .keyStatus_20_valid    (debounce_1_keyStatus_20_valid   ), //o
    .keyStatus_20_payload  (debounce_1_keyStatus_20_payload ), //o
    .keyStatus_21_valid    (debounce_1_keyStatus_21_valid   ), //o
    .keyStatus_21_payload  (debounce_1_keyStatus_21_payload ), //o
    .keyStatus_22_valid    (debounce_1_keyStatus_22_valid   ), //o
    .keyStatus_22_payload  (debounce_1_keyStatus_22_payload ), //o
    .keyStatus_23_valid    (debounce_1_keyStatus_23_valid   ), //o
    .keyStatus_23_payload  (debounce_1_keyStatus_23_payload ), //o
    .keyStatus_24_valid    (debounce_1_keyStatus_24_valid   ), //o
    .keyStatus_24_payload  (debounce_1_keyStatus_24_payload ), //o
    .keyStatus_25_valid    (debounce_1_keyStatus_25_valid   ), //o
    .keyStatus_25_payload  (debounce_1_keyStatus_25_payload ), //o
    .keyStatus_26_valid    (debounce_1_keyStatus_26_valid   ), //o
    .keyStatus_26_payload  (debounce_1_keyStatus_26_payload ), //o
    .keyStatus_27_valid    (debounce_1_keyStatus_27_valid   ), //o
    .keyStatus_27_payload  (debounce_1_keyStatus_27_payload ), //o
    .keyStatus_28_valid    (debounce_1_keyStatus_28_valid   ), //o
    .keyStatus_28_payload  (debounce_1_keyStatus_28_payload ), //o
    .keyStatus_29_valid    (debounce_1_keyStatus_29_valid   ), //o
    .keyStatus_29_payload  (debounce_1_keyStatus_29_payload ), //o
    .keyStatus_30_valid    (debounce_1_keyStatus_30_valid   ), //o
    .keyStatus_30_payload  (debounce_1_keyStatus_30_payload ), //o
    .keyStatus_31_valid    (debounce_1_keyStatus_31_valid   ), //o
    .keyStatus_31_payload  (debounce_1_keyStatus_31_payload ), //o
    .keyStatus_32_valid    (debounce_1_keyStatus_32_valid   ), //o
    .keyStatus_32_payload  (debounce_1_keyStatus_32_payload ), //o
    .keyStatus_33_valid    (debounce_1_keyStatus_33_valid   ), //o
    .keyStatus_33_payload  (debounce_1_keyStatus_33_payload ), //o
    .keyStatus_34_valid    (debounce_1_keyStatus_34_valid   ), //o
    .keyStatus_34_payload  (debounce_1_keyStatus_34_payload ), //o
    .keyStatus_35_valid    (debounce_1_keyStatus_35_valid   ), //o
    .keyStatus_35_payload  (debounce_1_keyStatus_35_payload ), //o
    .keyStatus_36_valid    (debounce_1_keyStatus_36_valid   ), //o
    .keyStatus_36_payload  (debounce_1_keyStatus_36_payload ), //o
    .keyStatus_37_valid    (debounce_1_keyStatus_37_valid   ), //o
    .keyStatus_37_payload  (debounce_1_keyStatus_37_payload ), //o
    .keyStatus_38_valid    (debounce_1_keyStatus_38_valid   ), //o
    .keyStatus_38_payload  (debounce_1_keyStatus_38_payload ), //o
    .keyStatus_39_valid    (debounce_1_keyStatus_39_valid   ), //o
    .keyStatus_39_payload  (debounce_1_keyStatus_39_payload ), //o
    .keyStatus_40_valid    (debounce_1_keyStatus_40_valid   ), //o
    .keyStatus_40_payload  (debounce_1_keyStatus_40_payload ), //o
    .keyStatus_41_valid    (debounce_1_keyStatus_41_valid   ), //o
    .keyStatus_41_payload  (debounce_1_keyStatus_41_payload ), //o
    .keyStatus_42_valid    (debounce_1_keyStatus_42_valid   ), //o
    .keyStatus_42_payload  (debounce_1_keyStatus_42_payload ), //o
    .keyStatus_43_valid    (debounce_1_keyStatus_43_valid   ), //o
    .keyStatus_43_payload  (debounce_1_keyStatus_43_payload ), //o
    .keyStatus_44_valid    (debounce_1_keyStatus_44_valid   ), //o
    .keyStatus_44_payload  (debounce_1_keyStatus_44_payload ), //o
    .keyStatus_45_valid    (debounce_1_keyStatus_45_valid   ), //o
    .keyStatus_45_payload  (debounce_1_keyStatus_45_payload ), //o
    .keyStatus_46_valid    (debounce_1_keyStatus_46_valid   ), //o
    .keyStatus_46_payload  (debounce_1_keyStatus_46_payload ), //o
    .keyStatus_47_valid    (debounce_1_keyStatus_47_valid   ), //o
    .keyStatus_47_payload  (debounce_1_keyStatus_47_payload ), //o
    .keyStatus_48_valid    (debounce_1_keyStatus_48_valid   ), //o
    .keyStatus_48_payload  (debounce_1_keyStatus_48_payload ), //o
    .keyStatus_49_valid    (debounce_1_keyStatus_49_valid   ), //o
    .keyStatus_49_payload  (debounce_1_keyStatus_49_payload ), //o
    .keyStatus_50_valid    (debounce_1_keyStatus_50_valid   ), //o
    .keyStatus_50_payload  (debounce_1_keyStatus_50_payload ), //o
    .keyStatus_51_valid    (debounce_1_keyStatus_51_valid   ), //o
    .keyStatus_51_payload  (debounce_1_keyStatus_51_payload ), //o
    .keyStatus_52_valid    (debounce_1_keyStatus_52_valid   ), //o
    .keyStatus_52_payload  (debounce_1_keyStatus_52_payload ), //o
    .keyStatus_53_valid    (debounce_1_keyStatus_53_valid   ), //o
    .keyStatus_53_payload  (debounce_1_keyStatus_53_payload ), //o
    .keyStatus_54_valid    (debounce_1_keyStatus_54_valid   ), //o
    .keyStatus_54_payload  (debounce_1_keyStatus_54_payload ), //o
    .keyStatus_55_valid    (debounce_1_keyStatus_55_valid   ), //o
    .keyStatus_55_payload  (debounce_1_keyStatus_55_payload ), //o
    .keyStatus_56_valid    (debounce_1_keyStatus_56_valid   ), //o
    .keyStatus_56_payload  (debounce_1_keyStatus_56_payload ), //o
    .keyStatus_57_valid    (debounce_1_keyStatus_57_valid   ), //o
    .keyStatus_57_payload  (debounce_1_keyStatus_57_payload ), //o
    .keyStatus_58_valid    (debounce_1_keyStatus_58_valid   ), //o
    .keyStatus_58_payload  (debounce_1_keyStatus_58_payload ), //o
    .keyStatus_59_valid    (debounce_1_keyStatus_59_valid   ), //o
    .keyStatus_59_payload  (debounce_1_keyStatus_59_payload ), //o
    .keyStatus_60_valid    (debounce_1_keyStatus_60_valid   ), //o
    .keyStatus_60_payload  (debounce_1_keyStatus_60_payload ), //o
    .keyStatus_61_valid    (debounce_1_keyStatus_61_valid   ), //o
    .keyStatus_61_payload  (debounce_1_keyStatus_61_payload ), //o
    .keyStatus_62_valid    (debounce_1_keyStatus_62_valid   ), //o
    .keyStatus_62_payload  (debounce_1_keyStatus_62_payload ), //o
    .keyStatus_63_valid    (debounce_1_keyStatus_63_valid   ), //o
    .keyStatus_63_payload  (debounce_1_keyStatus_63_payload ), //o
    .keyStatus_64_valid    (debounce_1_keyStatus_64_valid   ), //o
    .keyStatus_64_payload  (debounce_1_keyStatus_64_payload ), //o
    .keyStatus_65_valid    (debounce_1_keyStatus_65_valid   ), //o
    .keyStatus_65_payload  (debounce_1_keyStatus_65_payload ), //o
    .keyStatus_66_valid    (debounce_1_keyStatus_66_valid   ), //o
    .keyStatus_66_payload  (debounce_1_keyStatus_66_payload ), //o
    .keyStatus_67_valid    (debounce_1_keyStatus_67_valid   ), //o
    .keyStatus_67_payload  (debounce_1_keyStatus_67_payload ), //o
    .keyStatus_68_valid    (debounce_1_keyStatus_68_valid   ), //o
    .keyStatus_68_payload  (debounce_1_keyStatus_68_payload ), //o
    .keyStatus_69_valid    (debounce_1_keyStatus_69_valid   ), //o
    .keyStatus_69_payload  (debounce_1_keyStatus_69_payload ), //o
    .keyStatus_70_valid    (debounce_1_keyStatus_70_valid   ), //o
    .keyStatus_70_payload  (debounce_1_keyStatus_70_payload ), //o
    .keyStatus_71_valid    (debounce_1_keyStatus_71_valid   ), //o
    .keyStatus_71_payload  (debounce_1_keyStatus_71_payload ), //o
    .keyStatus_72_valid    (debounce_1_keyStatus_72_valid   ), //o
    .keyStatus_72_payload  (debounce_1_keyStatus_72_payload ), //o
    .keyStatus_73_valid    (debounce_1_keyStatus_73_valid   ), //o
    .keyStatus_73_payload  (debounce_1_keyStatus_73_payload ), //o
    .keyStatus_74_valid    (debounce_1_keyStatus_74_valid   ), //o
    .keyStatus_74_payload  (debounce_1_keyStatus_74_payload ), //o
    .keyStatus_75_valid    (debounce_1_keyStatus_75_valid   ), //o
    .keyStatus_75_payload  (debounce_1_keyStatus_75_payload ), //o
    .keyStatus_76_valid    (debounce_1_keyStatus_76_valid   ), //o
    .keyStatus_76_payload  (debounce_1_keyStatus_76_payload ), //o
    .keyStatus_77_valid    (debounce_1_keyStatus_77_valid   ), //o
    .keyStatus_77_payload  (debounce_1_keyStatus_77_payload ), //o
    .keyStatus_78_valid    (debounce_1_keyStatus_78_valid   ), //o
    .keyStatus_78_payload  (debounce_1_keyStatus_78_payload ), //o
    .keyStatus_79_valid    (debounce_1_keyStatus_79_valid   ), //o
    .keyStatus_79_payload  (debounce_1_keyStatus_79_payload ), //o
    .keyStatus_80_valid    (debounce_1_keyStatus_80_valid   ), //o
    .keyStatus_80_payload  (debounce_1_keyStatus_80_payload ), //o
    .keyStatus_81_valid    (debounce_1_keyStatus_81_valid   ), //o
    .keyStatus_81_payload  (debounce_1_keyStatus_81_payload ), //o
    .keyStatus_82_valid    (debounce_1_keyStatus_82_valid   ), //o
    .keyStatus_82_payload  (debounce_1_keyStatus_82_payload ), //o
    .keyStatus_83_valid    (debounce_1_keyStatus_83_valid   ), //o
    .keyStatus_83_payload  (debounce_1_keyStatus_83_payload ), //o
    .keyStatus_84_valid    (debounce_1_keyStatus_84_valid   ), //o
    .keyStatus_84_payload  (debounce_1_keyStatus_84_payload ), //o
    .keyStatus_85_valid    (debounce_1_keyStatus_85_valid   ), //o
    .keyStatus_85_payload  (debounce_1_keyStatus_85_payload ), //o
    .keyStatus_86_valid    (debounce_1_keyStatus_86_valid   ), //o
    .keyStatus_86_payload  (debounce_1_keyStatus_86_payload ), //o
    .keyStatus_87_valid    (debounce_1_keyStatus_87_valid   ), //o
    .keyStatus_87_payload  (debounce_1_keyStatus_87_payload ), //o
    .keyStatus_88_valid    (debounce_1_keyStatus_88_valid   ), //o
    .keyStatus_88_payload  (debounce_1_keyStatus_88_payload ), //o
    .keyStatus_89_valid    (debounce_1_keyStatus_89_valid   ), //o
    .keyStatus_89_payload  (debounce_1_keyStatus_89_payload ), //o
    .keyStatus_90_valid    (debounce_1_keyStatus_90_valid   ), //o
    .keyStatus_90_payload  (debounce_1_keyStatus_90_payload ), //o
    .keyStatus_91_valid    (debounce_1_keyStatus_91_valid   ), //o
    .keyStatus_91_payload  (debounce_1_keyStatus_91_payload ), //o
    .keyStatus_92_valid    (debounce_1_keyStatus_92_valid   ), //o
    .keyStatus_92_payload  (debounce_1_keyStatus_92_payload ), //o
    .keyStatus_93_valid    (debounce_1_keyStatus_93_valid   ), //o
    .keyStatus_93_payload  (debounce_1_keyStatus_93_payload ), //o
    .keyStatus_94_valid    (debounce_1_keyStatus_94_valid   ), //o
    .keyStatus_94_payload  (debounce_1_keyStatus_94_payload ), //o
    .keyStatus_95_valid    (debounce_1_keyStatus_95_valid   ), //o
    .keyStatus_95_payload  (debounce_1_keyStatus_95_payload ), //o
    .keyStatus_96_valid    (debounce_1_keyStatus_96_valid   ), //o
    .keyStatus_96_payload  (debounce_1_keyStatus_96_payload ), //o
    .keyStatus_97_valid    (debounce_1_keyStatus_97_valid   ), //o
    .keyStatus_97_payload  (debounce_1_keyStatus_97_payload ), //o
    .keyStatus_98_valid    (debounce_1_keyStatus_98_valid   ), //o
    .keyStatus_98_payload  (debounce_1_keyStatus_98_payload ), //o
    .keyStatus_99_valid    (debounce_1_keyStatus_99_valid   ), //o
    .keyStatus_99_payload  (debounce_1_keyStatus_99_payload ), //o
    .keyStatus_100_valid   (debounce_1_keyStatus_100_valid  ), //o
    .keyStatus_100_payload (debounce_1_keyStatus_100_payload), //o
    .keyStatus_101_valid   (debounce_1_keyStatus_101_valid  ), //o
    .keyStatus_101_payload (debounce_1_keyStatus_101_payload), //o
    .keyStatus_102_valid   (debounce_1_keyStatus_102_valid  ), //o
    .keyStatus_102_payload (debounce_1_keyStatus_102_payload), //o
    .CLK_50                (CLK_50                          ), //i
    ._zz_LED_R6            (_zz_LED_R6                      )  //i
  );
  always @(*) begin
    case(_zz_scanIdx_valid_2)
      7'b0000000 : begin
        _zz_scanIdx_valid_3 = keyStatus_0_valid;
        _zz_scanIdx_payload = keyStatus_0_payload;
      end
      7'b0000001 : begin
        _zz_scanIdx_valid_3 = keyStatus_1_valid;
        _zz_scanIdx_payload = keyStatus_1_payload;
      end
      7'b0000010 : begin
        _zz_scanIdx_valid_3 = keyStatus_2_valid;
        _zz_scanIdx_payload = keyStatus_2_payload;
      end
      7'b0000011 : begin
        _zz_scanIdx_valid_3 = keyStatus_3_valid;
        _zz_scanIdx_payload = keyStatus_3_payload;
      end
      7'b0000100 : begin
        _zz_scanIdx_valid_3 = keyStatus_4_valid;
        _zz_scanIdx_payload = keyStatus_4_payload;
      end
      7'b0000101 : begin
        _zz_scanIdx_valid_3 = keyStatus_5_valid;
        _zz_scanIdx_payload = keyStatus_5_payload;
      end
      7'b0000110 : begin
        _zz_scanIdx_valid_3 = keyStatus_6_valid;
        _zz_scanIdx_payload = keyStatus_6_payload;
      end
      7'b0000111 : begin
        _zz_scanIdx_valid_3 = keyStatus_7_valid;
        _zz_scanIdx_payload = keyStatus_7_payload;
      end
      7'b0001000 : begin
        _zz_scanIdx_valid_3 = keyStatus_8_valid;
        _zz_scanIdx_payload = keyStatus_8_payload;
      end
      7'b0001001 : begin
        _zz_scanIdx_valid_3 = keyStatus_9_valid;
        _zz_scanIdx_payload = keyStatus_9_payload;
      end
      7'b0001010 : begin
        _zz_scanIdx_valid_3 = keyStatus_10_valid;
        _zz_scanIdx_payload = keyStatus_10_payload;
      end
      7'b0001011 : begin
        _zz_scanIdx_valid_3 = keyStatus_11_valid;
        _zz_scanIdx_payload = keyStatus_11_payload;
      end
      7'b0001100 : begin
        _zz_scanIdx_valid_3 = keyStatus_12_valid;
        _zz_scanIdx_payload = keyStatus_12_payload;
      end
      7'b0001101 : begin
        _zz_scanIdx_valid_3 = keyStatus_13_valid;
        _zz_scanIdx_payload = keyStatus_13_payload;
      end
      7'b0001110 : begin
        _zz_scanIdx_valid_3 = keyStatus_14_valid;
        _zz_scanIdx_payload = keyStatus_14_payload;
      end
      7'b0001111 : begin
        _zz_scanIdx_valid_3 = keyStatus_15_valid;
        _zz_scanIdx_payload = keyStatus_15_payload;
      end
      7'b0010000 : begin
        _zz_scanIdx_valid_3 = keyStatus_16_valid;
        _zz_scanIdx_payload = keyStatus_16_payload;
      end
      7'b0010001 : begin
        _zz_scanIdx_valid_3 = keyStatus_17_valid;
        _zz_scanIdx_payload = keyStatus_17_payload;
      end
      7'b0010010 : begin
        _zz_scanIdx_valid_3 = keyStatus_18_valid;
        _zz_scanIdx_payload = keyStatus_18_payload;
      end
      7'b0010011 : begin
        _zz_scanIdx_valid_3 = keyStatus_19_valid;
        _zz_scanIdx_payload = keyStatus_19_payload;
      end
      7'b0010100 : begin
        _zz_scanIdx_valid_3 = keyStatus_20_valid;
        _zz_scanIdx_payload = keyStatus_20_payload;
      end
      7'b0010101 : begin
        _zz_scanIdx_valid_3 = keyStatus_21_valid;
        _zz_scanIdx_payload = keyStatus_21_payload;
      end
      7'b0010110 : begin
        _zz_scanIdx_valid_3 = keyStatus_22_valid;
        _zz_scanIdx_payload = keyStatus_22_payload;
      end
      7'b0010111 : begin
        _zz_scanIdx_valid_3 = keyStatus_23_valid;
        _zz_scanIdx_payload = keyStatus_23_payload;
      end
      7'b0011000 : begin
        _zz_scanIdx_valid_3 = keyStatus_24_valid;
        _zz_scanIdx_payload = keyStatus_24_payload;
      end
      7'b0011001 : begin
        _zz_scanIdx_valid_3 = keyStatus_25_valid;
        _zz_scanIdx_payload = keyStatus_25_payload;
      end
      7'b0011010 : begin
        _zz_scanIdx_valid_3 = keyStatus_26_valid;
        _zz_scanIdx_payload = keyStatus_26_payload;
      end
      7'b0011011 : begin
        _zz_scanIdx_valid_3 = keyStatus_27_valid;
        _zz_scanIdx_payload = keyStatus_27_payload;
      end
      7'b0011100 : begin
        _zz_scanIdx_valid_3 = keyStatus_28_valid;
        _zz_scanIdx_payload = keyStatus_28_payload;
      end
      7'b0011101 : begin
        _zz_scanIdx_valid_3 = keyStatus_29_valid;
        _zz_scanIdx_payload = keyStatus_29_payload;
      end
      7'b0011110 : begin
        _zz_scanIdx_valid_3 = keyStatus_30_valid;
        _zz_scanIdx_payload = keyStatus_30_payload;
      end
      7'b0011111 : begin
        _zz_scanIdx_valid_3 = keyStatus_31_valid;
        _zz_scanIdx_payload = keyStatus_31_payload;
      end
      7'b0100000 : begin
        _zz_scanIdx_valid_3 = keyStatus_32_valid;
        _zz_scanIdx_payload = keyStatus_32_payload;
      end
      7'b0100001 : begin
        _zz_scanIdx_valid_3 = keyStatus_33_valid;
        _zz_scanIdx_payload = keyStatus_33_payload;
      end
      7'b0100010 : begin
        _zz_scanIdx_valid_3 = keyStatus_34_valid;
        _zz_scanIdx_payload = keyStatus_34_payload;
      end
      7'b0100011 : begin
        _zz_scanIdx_valid_3 = keyStatus_35_valid;
        _zz_scanIdx_payload = keyStatus_35_payload;
      end
      7'b0100100 : begin
        _zz_scanIdx_valid_3 = keyStatus_36_valid;
        _zz_scanIdx_payload = keyStatus_36_payload;
      end
      7'b0100101 : begin
        _zz_scanIdx_valid_3 = keyStatus_37_valid;
        _zz_scanIdx_payload = keyStatus_37_payload;
      end
      7'b0100110 : begin
        _zz_scanIdx_valid_3 = keyStatus_38_valid;
        _zz_scanIdx_payload = keyStatus_38_payload;
      end
      7'b0100111 : begin
        _zz_scanIdx_valid_3 = keyStatus_39_valid;
        _zz_scanIdx_payload = keyStatus_39_payload;
      end
      7'b0101000 : begin
        _zz_scanIdx_valid_3 = keyStatus_40_valid;
        _zz_scanIdx_payload = keyStatus_40_payload;
      end
      7'b0101001 : begin
        _zz_scanIdx_valid_3 = keyStatus_41_valid;
        _zz_scanIdx_payload = keyStatus_41_payload;
      end
      7'b0101010 : begin
        _zz_scanIdx_valid_3 = keyStatus_42_valid;
        _zz_scanIdx_payload = keyStatus_42_payload;
      end
      7'b0101011 : begin
        _zz_scanIdx_valid_3 = keyStatus_43_valid;
        _zz_scanIdx_payload = keyStatus_43_payload;
      end
      7'b0101100 : begin
        _zz_scanIdx_valid_3 = keyStatus_44_valid;
        _zz_scanIdx_payload = keyStatus_44_payload;
      end
      7'b0101101 : begin
        _zz_scanIdx_valid_3 = keyStatus_45_valid;
        _zz_scanIdx_payload = keyStatus_45_payload;
      end
      7'b0101110 : begin
        _zz_scanIdx_valid_3 = keyStatus_46_valid;
        _zz_scanIdx_payload = keyStatus_46_payload;
      end
      7'b0101111 : begin
        _zz_scanIdx_valid_3 = keyStatus_47_valid;
        _zz_scanIdx_payload = keyStatus_47_payload;
      end
      7'b0110000 : begin
        _zz_scanIdx_valid_3 = keyStatus_48_valid;
        _zz_scanIdx_payload = keyStatus_48_payload;
      end
      7'b0110001 : begin
        _zz_scanIdx_valid_3 = keyStatus_49_valid;
        _zz_scanIdx_payload = keyStatus_49_payload;
      end
      7'b0110010 : begin
        _zz_scanIdx_valid_3 = keyStatus_50_valid;
        _zz_scanIdx_payload = keyStatus_50_payload;
      end
      7'b0110011 : begin
        _zz_scanIdx_valid_3 = keyStatus_51_valid;
        _zz_scanIdx_payload = keyStatus_51_payload;
      end
      7'b0110100 : begin
        _zz_scanIdx_valid_3 = keyStatus_52_valid;
        _zz_scanIdx_payload = keyStatus_52_payload;
      end
      7'b0110101 : begin
        _zz_scanIdx_valid_3 = keyStatus_53_valid;
        _zz_scanIdx_payload = keyStatus_53_payload;
      end
      7'b0110110 : begin
        _zz_scanIdx_valid_3 = keyStatus_54_valid;
        _zz_scanIdx_payload = keyStatus_54_payload;
      end
      7'b0110111 : begin
        _zz_scanIdx_valid_3 = keyStatus_55_valid;
        _zz_scanIdx_payload = keyStatus_55_payload;
      end
      7'b0111000 : begin
        _zz_scanIdx_valid_3 = keyStatus_56_valid;
        _zz_scanIdx_payload = keyStatus_56_payload;
      end
      7'b0111001 : begin
        _zz_scanIdx_valid_3 = keyStatus_57_valid;
        _zz_scanIdx_payload = keyStatus_57_payload;
      end
      7'b0111010 : begin
        _zz_scanIdx_valid_3 = keyStatus_58_valid;
        _zz_scanIdx_payload = keyStatus_58_payload;
      end
      7'b0111011 : begin
        _zz_scanIdx_valid_3 = keyStatus_59_valid;
        _zz_scanIdx_payload = keyStatus_59_payload;
      end
      7'b0111100 : begin
        _zz_scanIdx_valid_3 = keyStatus_60_valid;
        _zz_scanIdx_payload = keyStatus_60_payload;
      end
      7'b0111101 : begin
        _zz_scanIdx_valid_3 = keyStatus_61_valid;
        _zz_scanIdx_payload = keyStatus_61_payload;
      end
      7'b0111110 : begin
        _zz_scanIdx_valid_3 = keyStatus_62_valid;
        _zz_scanIdx_payload = keyStatus_62_payload;
      end
      7'b0111111 : begin
        _zz_scanIdx_valid_3 = keyStatus_63_valid;
        _zz_scanIdx_payload = keyStatus_63_payload;
      end
      7'b1000000 : begin
        _zz_scanIdx_valid_3 = keyStatus_64_valid;
        _zz_scanIdx_payload = keyStatus_64_payload;
      end
      7'b1000001 : begin
        _zz_scanIdx_valid_3 = keyStatus_65_valid;
        _zz_scanIdx_payload = keyStatus_65_payload;
      end
      7'b1000010 : begin
        _zz_scanIdx_valid_3 = keyStatus_66_valid;
        _zz_scanIdx_payload = keyStatus_66_payload;
      end
      7'b1000011 : begin
        _zz_scanIdx_valid_3 = keyStatus_67_valid;
        _zz_scanIdx_payload = keyStatus_67_payload;
      end
      7'b1000100 : begin
        _zz_scanIdx_valid_3 = keyStatus_68_valid;
        _zz_scanIdx_payload = keyStatus_68_payload;
      end
      7'b1000101 : begin
        _zz_scanIdx_valid_3 = keyStatus_69_valid;
        _zz_scanIdx_payload = keyStatus_69_payload;
      end
      7'b1000110 : begin
        _zz_scanIdx_valid_3 = keyStatus_70_valid;
        _zz_scanIdx_payload = keyStatus_70_payload;
      end
      7'b1000111 : begin
        _zz_scanIdx_valid_3 = keyStatus_71_valid;
        _zz_scanIdx_payload = keyStatus_71_payload;
      end
      7'b1001000 : begin
        _zz_scanIdx_valid_3 = keyStatus_72_valid;
        _zz_scanIdx_payload = keyStatus_72_payload;
      end
      7'b1001001 : begin
        _zz_scanIdx_valid_3 = keyStatus_73_valid;
        _zz_scanIdx_payload = keyStatus_73_payload;
      end
      7'b1001010 : begin
        _zz_scanIdx_valid_3 = keyStatus_74_valid;
        _zz_scanIdx_payload = keyStatus_74_payload;
      end
      7'b1001011 : begin
        _zz_scanIdx_valid_3 = keyStatus_75_valid;
        _zz_scanIdx_payload = keyStatus_75_payload;
      end
      7'b1001100 : begin
        _zz_scanIdx_valid_3 = keyStatus_76_valid;
        _zz_scanIdx_payload = keyStatus_76_payload;
      end
      7'b1001101 : begin
        _zz_scanIdx_valid_3 = keyStatus_77_valid;
        _zz_scanIdx_payload = keyStatus_77_payload;
      end
      7'b1001110 : begin
        _zz_scanIdx_valid_3 = keyStatus_78_valid;
        _zz_scanIdx_payload = keyStatus_78_payload;
      end
      7'b1001111 : begin
        _zz_scanIdx_valid_3 = keyStatus_79_valid;
        _zz_scanIdx_payload = keyStatus_79_payload;
      end
      7'b1010000 : begin
        _zz_scanIdx_valid_3 = keyStatus_80_valid;
        _zz_scanIdx_payload = keyStatus_80_payload;
      end
      7'b1010001 : begin
        _zz_scanIdx_valid_3 = keyStatus_81_valid;
        _zz_scanIdx_payload = keyStatus_81_payload;
      end
      7'b1010010 : begin
        _zz_scanIdx_valid_3 = keyStatus_82_valid;
        _zz_scanIdx_payload = keyStatus_82_payload;
      end
      7'b1010011 : begin
        _zz_scanIdx_valid_3 = keyStatus_83_valid;
        _zz_scanIdx_payload = keyStatus_83_payload;
      end
      7'b1010100 : begin
        _zz_scanIdx_valid_3 = keyStatus_84_valid;
        _zz_scanIdx_payload = keyStatus_84_payload;
      end
      7'b1010101 : begin
        _zz_scanIdx_valid_3 = keyStatus_85_valid;
        _zz_scanIdx_payload = keyStatus_85_payload;
      end
      7'b1010110 : begin
        _zz_scanIdx_valid_3 = keyStatus_86_valid;
        _zz_scanIdx_payload = keyStatus_86_payload;
      end
      7'b1010111 : begin
        _zz_scanIdx_valid_3 = keyStatus_87_valid;
        _zz_scanIdx_payload = keyStatus_87_payload;
      end
      7'b1011000 : begin
        _zz_scanIdx_valid_3 = keyStatus_88_valid;
        _zz_scanIdx_payload = keyStatus_88_payload;
      end
      7'b1011001 : begin
        _zz_scanIdx_valid_3 = keyStatus_89_valid;
        _zz_scanIdx_payload = keyStatus_89_payload;
      end
      7'b1011010 : begin
        _zz_scanIdx_valid_3 = keyStatus_90_valid;
        _zz_scanIdx_payload = keyStatus_90_payload;
      end
      7'b1011011 : begin
        _zz_scanIdx_valid_3 = keyStatus_91_valid;
        _zz_scanIdx_payload = keyStatus_91_payload;
      end
      7'b1011100 : begin
        _zz_scanIdx_valid_3 = keyStatus_92_valid;
        _zz_scanIdx_payload = keyStatus_92_payload;
      end
      7'b1011101 : begin
        _zz_scanIdx_valid_3 = keyStatus_93_valid;
        _zz_scanIdx_payload = keyStatus_93_payload;
      end
      7'b1011110 : begin
        _zz_scanIdx_valid_3 = keyStatus_94_valid;
        _zz_scanIdx_payload = keyStatus_94_payload;
      end
      7'b1011111 : begin
        _zz_scanIdx_valid_3 = keyStatus_95_valid;
        _zz_scanIdx_payload = keyStatus_95_payload;
      end
      7'b1100000 : begin
        _zz_scanIdx_valid_3 = keyStatus_96_valid;
        _zz_scanIdx_payload = keyStatus_96_payload;
      end
      7'b1100001 : begin
        _zz_scanIdx_valid_3 = keyStatus_97_valid;
        _zz_scanIdx_payload = keyStatus_97_payload;
      end
      7'b1100010 : begin
        _zz_scanIdx_valid_3 = keyStatus_98_valid;
        _zz_scanIdx_payload = keyStatus_98_payload;
      end
      7'b1100011 : begin
        _zz_scanIdx_valid_3 = keyStatus_99_valid;
        _zz_scanIdx_payload = keyStatus_99_payload;
      end
      7'b1100100 : begin
        _zz_scanIdx_valid_3 = keyStatus_100_valid;
        _zz_scanIdx_payload = keyStatus_100_payload;
      end
      7'b1100101 : begin
        _zz_scanIdx_valid_3 = keyStatus_101_valid;
        _zz_scanIdx_payload = keyStatus_101_payload;
      end
      default : begin
        _zz_scanIdx_valid_3 = keyStatus_102_valid;
        _zz_scanIdx_payload = keyStatus_102_payload;
      end
    endcase
  end

  always @(*) begin
    clkScan_stateRise = 1'b0;
    if(clkScan_counter_willOverflow) begin
      clkScan_stateRise = (! clkScan_state);
    end
    if(clkScan_state) begin
      clkScan_stateRise = 1'b0;
    end
  end

  always @(*) begin
    clkScan_counter_willClear = 1'b0;
    if(clkScan_state) begin
      clkScan_counter_willClear = 1'b1;
    end
  end

  assign clkScan_counter_willOverflowIfInc = (clkScan_counter_value == 13'h1045);
  assign clkScan_counter_willOverflow = (clkScan_counter_willOverflowIfInc && clkScan_counter_willIncrement);
  always @(*) begin
    if(clkScan_counter_willOverflow) begin
      clkScan_counter_valueNext = 13'h0;
    end else begin
      clkScan_counter_valueNext = (clkScan_counter_value + _zz_clkScan_counter_valueNext);
    end
    if(clkScan_counter_willClear) begin
      clkScan_counter_valueNext = 13'h0;
    end
  end

  assign clkScan_counter_willIncrement = 1'b1;
  assign ROW = scanK_ROW;
  assign keyStatus_0_valid = debounce_1_keyStatus_0_valid;
  assign keyStatus_0_payload = debounce_1_keyStatus_0_payload;
  assign keyStatus_1_valid = debounce_1_keyStatus_1_valid;
  assign keyStatus_1_payload = debounce_1_keyStatus_1_payload;
  assign keyStatus_2_valid = debounce_1_keyStatus_2_valid;
  assign keyStatus_2_payload = debounce_1_keyStatus_2_payload;
  assign keyStatus_3_valid = debounce_1_keyStatus_3_valid;
  assign keyStatus_3_payload = debounce_1_keyStatus_3_payload;
  assign keyStatus_4_valid = debounce_1_keyStatus_4_valid;
  assign keyStatus_4_payload = debounce_1_keyStatus_4_payload;
  assign keyStatus_5_valid = debounce_1_keyStatus_5_valid;
  assign keyStatus_5_payload = debounce_1_keyStatus_5_payload;
  assign keyStatus_6_valid = debounce_1_keyStatus_6_valid;
  assign keyStatus_6_payload = debounce_1_keyStatus_6_payload;
  assign keyStatus_7_valid = debounce_1_keyStatus_7_valid;
  assign keyStatus_7_payload = debounce_1_keyStatus_7_payload;
  assign keyStatus_8_valid = debounce_1_keyStatus_8_valid;
  assign keyStatus_8_payload = debounce_1_keyStatus_8_payload;
  assign keyStatus_9_valid = debounce_1_keyStatus_9_valid;
  assign keyStatus_9_payload = debounce_1_keyStatus_9_payload;
  assign keyStatus_10_valid = debounce_1_keyStatus_10_valid;
  assign keyStatus_10_payload = debounce_1_keyStatus_10_payload;
  assign keyStatus_11_valid = debounce_1_keyStatus_11_valid;
  assign keyStatus_11_payload = debounce_1_keyStatus_11_payload;
  assign keyStatus_12_valid = debounce_1_keyStatus_12_valid;
  assign keyStatus_12_payload = debounce_1_keyStatus_12_payload;
  assign keyStatus_13_valid = debounce_1_keyStatus_13_valid;
  assign keyStatus_13_payload = debounce_1_keyStatus_13_payload;
  assign keyStatus_14_valid = debounce_1_keyStatus_14_valid;
  assign keyStatus_14_payload = debounce_1_keyStatus_14_payload;
  assign keyStatus_15_valid = debounce_1_keyStatus_15_valid;
  assign keyStatus_15_payload = debounce_1_keyStatus_15_payload;
  assign keyStatus_16_valid = debounce_1_keyStatus_16_valid;
  assign keyStatus_16_payload = debounce_1_keyStatus_16_payload;
  assign keyStatus_17_valid = debounce_1_keyStatus_17_valid;
  assign keyStatus_17_payload = debounce_1_keyStatus_17_payload;
  assign keyStatus_18_valid = debounce_1_keyStatus_18_valid;
  assign keyStatus_18_payload = debounce_1_keyStatus_18_payload;
  assign keyStatus_19_valid = debounce_1_keyStatus_19_valid;
  assign keyStatus_19_payload = debounce_1_keyStatus_19_payload;
  assign keyStatus_20_valid = debounce_1_keyStatus_20_valid;
  assign keyStatus_20_payload = debounce_1_keyStatus_20_payload;
  assign keyStatus_21_valid = debounce_1_keyStatus_21_valid;
  assign keyStatus_21_payload = debounce_1_keyStatus_21_payload;
  assign keyStatus_22_valid = debounce_1_keyStatus_22_valid;
  assign keyStatus_22_payload = debounce_1_keyStatus_22_payload;
  assign keyStatus_23_valid = debounce_1_keyStatus_23_valid;
  assign keyStatus_23_payload = debounce_1_keyStatus_23_payload;
  assign keyStatus_24_valid = debounce_1_keyStatus_24_valid;
  assign keyStatus_24_payload = debounce_1_keyStatus_24_payload;
  assign keyStatus_25_valid = debounce_1_keyStatus_25_valid;
  assign keyStatus_25_payload = debounce_1_keyStatus_25_payload;
  assign keyStatus_26_valid = debounce_1_keyStatus_26_valid;
  assign keyStatus_26_payload = debounce_1_keyStatus_26_payload;
  assign keyStatus_27_valid = debounce_1_keyStatus_27_valid;
  assign keyStatus_27_payload = debounce_1_keyStatus_27_payload;
  assign keyStatus_28_valid = debounce_1_keyStatus_28_valid;
  assign keyStatus_28_payload = debounce_1_keyStatus_28_payload;
  assign keyStatus_29_valid = debounce_1_keyStatus_29_valid;
  assign keyStatus_29_payload = debounce_1_keyStatus_29_payload;
  assign keyStatus_30_valid = debounce_1_keyStatus_30_valid;
  assign keyStatus_30_payload = debounce_1_keyStatus_30_payload;
  assign keyStatus_31_valid = debounce_1_keyStatus_31_valid;
  assign keyStatus_31_payload = debounce_1_keyStatus_31_payload;
  assign keyStatus_32_valid = debounce_1_keyStatus_32_valid;
  assign keyStatus_32_payload = debounce_1_keyStatus_32_payload;
  assign keyStatus_33_valid = debounce_1_keyStatus_33_valid;
  assign keyStatus_33_payload = debounce_1_keyStatus_33_payload;
  assign keyStatus_34_valid = debounce_1_keyStatus_34_valid;
  assign keyStatus_34_payload = debounce_1_keyStatus_34_payload;
  assign keyStatus_35_valid = debounce_1_keyStatus_35_valid;
  assign keyStatus_35_payload = debounce_1_keyStatus_35_payload;
  assign keyStatus_36_valid = debounce_1_keyStatus_36_valid;
  assign keyStatus_36_payload = debounce_1_keyStatus_36_payload;
  assign keyStatus_37_valid = debounce_1_keyStatus_37_valid;
  assign keyStatus_37_payload = debounce_1_keyStatus_37_payload;
  assign keyStatus_38_valid = debounce_1_keyStatus_38_valid;
  assign keyStatus_38_payload = debounce_1_keyStatus_38_payload;
  assign keyStatus_39_valid = debounce_1_keyStatus_39_valid;
  assign keyStatus_39_payload = debounce_1_keyStatus_39_payload;
  assign keyStatus_40_valid = debounce_1_keyStatus_40_valid;
  assign keyStatus_40_payload = debounce_1_keyStatus_40_payload;
  assign keyStatus_41_valid = debounce_1_keyStatus_41_valid;
  assign keyStatus_41_payload = debounce_1_keyStatus_41_payload;
  assign keyStatus_42_valid = debounce_1_keyStatus_42_valid;
  assign keyStatus_42_payload = debounce_1_keyStatus_42_payload;
  assign keyStatus_43_valid = debounce_1_keyStatus_43_valid;
  assign keyStatus_43_payload = debounce_1_keyStatus_43_payload;
  assign keyStatus_44_valid = debounce_1_keyStatus_44_valid;
  assign keyStatus_44_payload = debounce_1_keyStatus_44_payload;
  assign keyStatus_45_valid = debounce_1_keyStatus_45_valid;
  assign keyStatus_45_payload = debounce_1_keyStatus_45_payload;
  assign keyStatus_46_valid = debounce_1_keyStatus_46_valid;
  assign keyStatus_46_payload = debounce_1_keyStatus_46_payload;
  assign keyStatus_47_valid = debounce_1_keyStatus_47_valid;
  assign keyStatus_47_payload = debounce_1_keyStatus_47_payload;
  assign keyStatus_48_valid = debounce_1_keyStatus_48_valid;
  assign keyStatus_48_payload = debounce_1_keyStatus_48_payload;
  assign keyStatus_49_valid = debounce_1_keyStatus_49_valid;
  assign keyStatus_49_payload = debounce_1_keyStatus_49_payload;
  assign keyStatus_50_valid = debounce_1_keyStatus_50_valid;
  assign keyStatus_50_payload = debounce_1_keyStatus_50_payload;
  assign keyStatus_51_valid = debounce_1_keyStatus_51_valid;
  assign keyStatus_51_payload = debounce_1_keyStatus_51_payload;
  assign keyStatus_52_valid = debounce_1_keyStatus_52_valid;
  assign keyStatus_52_payload = debounce_1_keyStatus_52_payload;
  assign keyStatus_53_valid = debounce_1_keyStatus_53_valid;
  assign keyStatus_53_payload = debounce_1_keyStatus_53_payload;
  assign keyStatus_54_valid = debounce_1_keyStatus_54_valid;
  assign keyStatus_54_payload = debounce_1_keyStatus_54_payload;
  assign keyStatus_55_valid = debounce_1_keyStatus_55_valid;
  assign keyStatus_55_payload = debounce_1_keyStatus_55_payload;
  assign keyStatus_56_valid = debounce_1_keyStatus_56_valid;
  assign keyStatus_56_payload = debounce_1_keyStatus_56_payload;
  assign keyStatus_57_valid = debounce_1_keyStatus_57_valid;
  assign keyStatus_57_payload = debounce_1_keyStatus_57_payload;
  assign keyStatus_58_valid = debounce_1_keyStatus_58_valid;
  assign keyStatus_58_payload = debounce_1_keyStatus_58_payload;
  assign keyStatus_59_valid = debounce_1_keyStatus_59_valid;
  assign keyStatus_59_payload = debounce_1_keyStatus_59_payload;
  assign keyStatus_60_valid = debounce_1_keyStatus_60_valid;
  assign keyStatus_60_payload = debounce_1_keyStatus_60_payload;
  assign keyStatus_61_valid = debounce_1_keyStatus_61_valid;
  assign keyStatus_61_payload = debounce_1_keyStatus_61_payload;
  assign keyStatus_62_valid = debounce_1_keyStatus_62_valid;
  assign keyStatus_62_payload = debounce_1_keyStatus_62_payload;
  assign keyStatus_63_valid = debounce_1_keyStatus_63_valid;
  assign keyStatus_63_payload = debounce_1_keyStatus_63_payload;
  assign keyStatus_64_valid = debounce_1_keyStatus_64_valid;
  assign keyStatus_64_payload = debounce_1_keyStatus_64_payload;
  assign keyStatus_65_valid = debounce_1_keyStatus_65_valid;
  assign keyStatus_65_payload = debounce_1_keyStatus_65_payload;
  assign keyStatus_66_valid = debounce_1_keyStatus_66_valid;
  assign keyStatus_66_payload = debounce_1_keyStatus_66_payload;
  assign keyStatus_67_valid = debounce_1_keyStatus_67_valid;
  assign keyStatus_67_payload = debounce_1_keyStatus_67_payload;
  assign keyStatus_68_valid = debounce_1_keyStatus_68_valid;
  assign keyStatus_68_payload = debounce_1_keyStatus_68_payload;
  assign keyStatus_69_valid = debounce_1_keyStatus_69_valid;
  assign keyStatus_69_payload = debounce_1_keyStatus_69_payload;
  assign keyStatus_70_valid = debounce_1_keyStatus_70_valid;
  assign keyStatus_70_payload = debounce_1_keyStatus_70_payload;
  assign keyStatus_71_valid = debounce_1_keyStatus_71_valid;
  assign keyStatus_71_payload = debounce_1_keyStatus_71_payload;
  assign keyStatus_72_valid = debounce_1_keyStatus_72_valid;
  assign keyStatus_72_payload = debounce_1_keyStatus_72_payload;
  assign keyStatus_73_valid = debounce_1_keyStatus_73_valid;
  assign keyStatus_73_payload = debounce_1_keyStatus_73_payload;
  assign keyStatus_74_valid = debounce_1_keyStatus_74_valid;
  assign keyStatus_74_payload = debounce_1_keyStatus_74_payload;
  assign keyStatus_75_valid = debounce_1_keyStatus_75_valid;
  assign keyStatus_75_payload = debounce_1_keyStatus_75_payload;
  assign keyStatus_76_valid = debounce_1_keyStatus_76_valid;
  assign keyStatus_76_payload = debounce_1_keyStatus_76_payload;
  assign keyStatus_77_valid = debounce_1_keyStatus_77_valid;
  assign keyStatus_77_payload = debounce_1_keyStatus_77_payload;
  assign keyStatus_78_valid = debounce_1_keyStatus_78_valid;
  assign keyStatus_78_payload = debounce_1_keyStatus_78_payload;
  assign keyStatus_79_valid = debounce_1_keyStatus_79_valid;
  assign keyStatus_79_payload = debounce_1_keyStatus_79_payload;
  assign keyStatus_80_valid = debounce_1_keyStatus_80_valid;
  assign keyStatus_80_payload = debounce_1_keyStatus_80_payload;
  assign keyStatus_81_valid = debounce_1_keyStatus_81_valid;
  assign keyStatus_81_payload = debounce_1_keyStatus_81_payload;
  assign keyStatus_82_valid = debounce_1_keyStatus_82_valid;
  assign keyStatus_82_payload = debounce_1_keyStatus_82_payload;
  assign keyStatus_83_valid = debounce_1_keyStatus_83_valid;
  assign keyStatus_83_payload = debounce_1_keyStatus_83_payload;
  assign keyStatus_84_valid = debounce_1_keyStatus_84_valid;
  assign keyStatus_84_payload = debounce_1_keyStatus_84_payload;
  assign keyStatus_85_valid = debounce_1_keyStatus_85_valid;
  assign keyStatus_85_payload = debounce_1_keyStatus_85_payload;
  assign keyStatus_86_valid = debounce_1_keyStatus_86_valid;
  assign keyStatus_86_payload = debounce_1_keyStatus_86_payload;
  assign keyStatus_87_valid = debounce_1_keyStatus_87_valid;
  assign keyStatus_87_payload = debounce_1_keyStatus_87_payload;
  assign keyStatus_88_valid = debounce_1_keyStatus_88_valid;
  assign keyStatus_88_payload = debounce_1_keyStatus_88_payload;
  assign keyStatus_89_valid = debounce_1_keyStatus_89_valid;
  assign keyStatus_89_payload = debounce_1_keyStatus_89_payload;
  assign keyStatus_90_valid = debounce_1_keyStatus_90_valid;
  assign keyStatus_90_payload = debounce_1_keyStatus_90_payload;
  assign keyStatus_91_valid = debounce_1_keyStatus_91_valid;
  assign keyStatus_91_payload = debounce_1_keyStatus_91_payload;
  assign keyStatus_92_valid = debounce_1_keyStatus_92_valid;
  assign keyStatus_92_payload = debounce_1_keyStatus_92_payload;
  assign keyStatus_93_valid = debounce_1_keyStatus_93_valid;
  assign keyStatus_93_payload = debounce_1_keyStatus_93_payload;
  assign keyStatus_94_valid = debounce_1_keyStatus_94_valid;
  assign keyStatus_94_payload = debounce_1_keyStatus_94_payload;
  assign keyStatus_95_valid = debounce_1_keyStatus_95_valid;
  assign keyStatus_95_payload = debounce_1_keyStatus_95_payload;
  assign keyStatus_96_valid = debounce_1_keyStatus_96_valid;
  assign keyStatus_96_payload = debounce_1_keyStatus_96_payload;
  assign keyStatus_97_valid = debounce_1_keyStatus_97_valid;
  assign keyStatus_97_payload = debounce_1_keyStatus_97_payload;
  assign keyStatus_98_valid = debounce_1_keyStatus_98_valid;
  assign keyStatus_98_payload = debounce_1_keyStatus_98_payload;
  assign keyStatus_99_valid = debounce_1_keyStatus_99_valid;
  assign keyStatus_99_payload = debounce_1_keyStatus_99_payload;
  assign keyStatus_100_valid = debounce_1_keyStatus_100_valid;
  assign keyStatus_100_payload = debounce_1_keyStatus_100_payload;
  assign keyStatus_101_valid = debounce_1_keyStatus_101_valid;
  assign keyStatus_101_payload = debounce_1_keyStatus_101_payload;
  assign keyStatus_102_valid = debounce_1_keyStatus_102_valid;
  assign keyStatus_102_payload = debounce_1_keyStatus_102_payload;
  assign when_ClockDomain_l369 = (_zz_when_ClockDomain_l369 == 8'hf1);
  assign _zz_1 = (_zz_scanIdx_valid_2 == 7'h66);
  assign _zz_2 = (_zz_1 && _zz_scanIdx_valid);
  always @(*) begin
    if(_zz_2) begin
      _zz_scanIdx_valid_1 = 7'h0;
    end else begin
      _zz_scanIdx_valid_1 = (_zz_scanIdx_valid_2 + _zz__zz_scanIdx_valid_1);
    end
    if(1'b0) begin
      _zz_scanIdx_valid_1 = 7'h0;
    end
  end

  assign _zz_scanIdx_valid = 1'b1;
  assign scanIdx_valid = _zz_scanIdx_valid_3;
  assign scanIdx_payload = {_zz_scanIdx_payload,_zz_scanIdx_valid_2};
  always @(posedge CLK_50 or posedge _zz_LED_R6) begin
    if(_zz_LED_R6) begin
      clkScan_state <= 1'b0;
      clkScan_counter_value <= 13'h0;
      _zz_when_ClockDomain_l369 <= 8'h0;
      when_ClockDomain_l369_regNext <= 1'b0;
    end else begin
      clkScan_counter_value <= clkScan_counter_valueNext;
      if(clkScan_counter_willOverflow) begin
        clkScan_state <= 1'b1;
      end
      if(clkScan_state) begin
        clkScan_state <= 1'b0;
      end
      _zz_when_ClockDomain_l369 <= (_zz_when_ClockDomain_l369 + 8'h01);
      if(when_ClockDomain_l369) begin
        _zz_when_ClockDomain_l369 <= 8'h0;
      end
      when_ClockDomain_l369_regNext <= when_ClockDomain_l369;
    end
  end

  always @(posedge CLK_50 or posedge _zz_LED_R6) begin
    if(_zz_LED_R6) begin
      _zz_scanIdx_valid_2 <= 7'h0;
    end else begin
      if(when_ClockDomain_l369_regNext) begin
        _zz_scanIdx_valid_2 <= _zz_scanIdx_valid_1;
      end
    end
  end


endmodule

module BufferCC (
  input               io_dataIn,
  output              io_dataOut,
  input               CLK_50,
  input               _zz_1
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge CLK_50 or posedge _zz_1) begin
    if(_zz_1) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module ResetController (
  input               io_clock,
  input               io_externalReset,
  output              io_globalReset
);

  wire       [15:0]   _zz__zz_2;
  wire       [0:0]    _zz__zz_2_1;
  wire       [27:0]   _zz__zz_io_globalReset_2;
  wire       [0:0]    _zz__zz_io_globalReset_2_1;
  reg                 _zz_1;
  reg        [15:0]   _zz_2;
  reg        [15:0]   _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  reg                 _zz_io_globalReset;
  reg                 _zz_io_globalReset_1;
  reg                 _zz_6;
  reg        [27:0]   _zz_io_globalReset_2;
  reg        [27:0]   _zz_io_globalReset_3;
  wire                _zz_io_globalReset_4;
  wire                _zz_io_globalReset_5;
  reg                 io_externalReset_regNext;
  wire                when_ResetController_l26;
  reg                 _zz_io_globalReset_6;

  assign _zz__zz_2_1 = _zz_1;
  assign _zz__zz_2 = {15'd0, _zz__zz_2_1};
  assign _zz__zz_io_globalReset_2_1 = _zz_io_globalReset_1;
  assign _zz__zz_io_globalReset_2 = {27'd0, _zz__zz_io_globalReset_2_1};
  initial begin
    _zz_3 = 16'h0;
    _zz_io_globalReset = 1'b1;
    _zz_io_globalReset_3 = 28'h0;
    io_externalReset_regNext = 1'b0;
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(_zz_io_globalReset) begin
      _zz_1 = 1'b1;
    end
  end

  assign _zz_4 = (_zz_3 == 16'hc34f);
  assign _zz_5 = (_zz_4 && _zz_1);
  always @(*) begin
    if(_zz_5) begin
      _zz_2 = 16'h0;
    end else begin
      _zz_2 = (_zz_3 + _zz__zz_2);
    end
    if(1'b0) begin
      _zz_2 = 16'h0;
    end
  end

  always @(*) begin
    _zz_io_globalReset_1 = 1'b0;
    if(io_externalReset) begin
      _zz_io_globalReset_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_6 = 1'b0;
    if(when_ResetController_l26) begin
      _zz_6 = 1'b1;
    end
  end

  assign _zz_io_globalReset_4 = (_zz_io_globalReset_3 == 28'h8f0d17f);
  assign _zz_io_globalReset_5 = (_zz_io_globalReset_4 && _zz_io_globalReset_1);
  always @(*) begin
    if(_zz_io_globalReset_5) begin
      _zz_io_globalReset_2 = 28'h0;
    end else begin
      _zz_io_globalReset_2 = (_zz_io_globalReset_3 + _zz__zz_io_globalReset_2);
    end
    if(_zz_6) begin
      _zz_io_globalReset_2 = 28'h0;
    end
  end

  assign when_ResetController_l26 = (io_externalReset && (! io_externalReset_regNext));
  assign io_globalReset = _zz_io_globalReset_6;
  always @(posedge io_clock) begin
    _zz_3 <= _zz_2;
    if(_zz_4) begin
      _zz_io_globalReset <= 1'b0;
    end
    _zz_io_globalReset_3 <= _zz_io_globalReset_2;
    io_externalReset_regNext <= io_externalReset;
  end

  always @(posedge io_clock) begin
    _zz_io_globalReset_6 <= (_zz_io_globalReset || _zz_io_globalReset_5);
  end


endmodule

module UartCtrl_1 (
  input      [2:0]    io_config_frame_dataLength,
  input      [0:0]    io_config_frame_stop,
  input      [1:0]    io_config_frame_parity,
  input      [19:0]   io_config_clockDivider,
  input               io_write_valid,
  output reg          io_write_ready,
  input      [7:0]    io_write_payload,
  output              io_read_valid,
  input               io_read_ready,
  output     [7:0]    io_read_payload,
  output              io_uart_txd,
  input               io_uart_rxd,
  output              io_readError,
  input               io_writeBreak,
  output              io_readBreak,
  input               CLK_50,
  input               _zz_LED_R6
);
  localparam UartStopType_ONE = 1'd0;
  localparam UartStopType_TWO = 1'd1;
  localparam UartParityType_NONE = 2'd0;
  localparam UartParityType_EVEN = 2'd1;
  localparam UartParityType_ODD = 2'd2;

  wire                tx_io_write_ready;
  wire                tx_io_txd;
  wire                rx_io_read_valid;
  wire       [7:0]    rx_io_read_payload;
  wire                rx_io_rts;
  wire                rx_io_error;
  wire                rx_io_break;
  reg        [19:0]   clockDivider_counter;
  wire                clockDivider_tick;
  reg                 clockDivider_tickReg;
  reg                 io_write_thrown_valid;
  wire                io_write_thrown_ready;
  wire       [7:0]    io_write_thrown_payload;
  `ifndef SYNTHESIS
  reg [23:0] io_config_frame_stop_string;
  reg [31:0] io_config_frame_parity_string;
  `endif


  UartCtrlTx_1 tx (
    .io_configFrame_dataLength (io_config_frame_dataLength[2:0]), //i
    .io_configFrame_stop       (io_config_frame_stop           ), //i
    .io_configFrame_parity     (io_config_frame_parity[1:0]    ), //i
    .io_samplingTick           (clockDivider_tickReg           ), //i
    .io_write_valid            (io_write_thrown_valid          ), //i
    .io_write_ready            (tx_io_write_ready              ), //o
    .io_write_payload          (io_write_thrown_payload[7:0]   ), //i
    .io_cts                    (1'b0                           ), //i
    .io_txd                    (tx_io_txd                      ), //o
    .io_break                  (io_writeBreak                  ), //i
    .CLK_50                    (CLK_50                         ), //i
    ._zz_LED_R6                (_zz_LED_R6                     )  //i
  );
  UartCtrlRx_1 rx (
    .io_configFrame_dataLength (io_config_frame_dataLength[2:0]), //i
    .io_configFrame_stop       (io_config_frame_stop           ), //i
    .io_configFrame_parity     (io_config_frame_parity[1:0]    ), //i
    .io_samplingTick           (clockDivider_tickReg           ), //i
    .io_read_valid             (rx_io_read_valid               ), //o
    .io_read_ready             (io_read_ready                  ), //i
    .io_read_payload           (rx_io_read_payload[7:0]        ), //o
    .io_rxd                    (io_uart_rxd                    ), //i
    .io_rts                    (rx_io_rts                      ), //o
    .io_error                  (rx_io_error                    ), //o
    .io_break                  (rx_io_break                    ), //o
    .CLK_50                    (CLK_50                         ), //i
    ._zz_LED_R6                (_zz_LED_R6                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_config_frame_stop)
      UartStopType_ONE : io_config_frame_stop_string = "ONE";
      UartStopType_TWO : io_config_frame_stop_string = "TWO";
      default : io_config_frame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_config_frame_parity)
      UartParityType_NONE : io_config_frame_parity_string = "NONE";
      UartParityType_EVEN : io_config_frame_parity_string = "EVEN";
      UartParityType_ODD : io_config_frame_parity_string = "ODD ";
      default : io_config_frame_parity_string = "????";
    endcase
  end
  `endif

  assign clockDivider_tick = (clockDivider_counter == 20'h0);
  always @(*) begin
    io_write_thrown_valid = io_write_valid;
    if(rx_io_break) begin
      io_write_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    io_write_ready = io_write_thrown_ready;
    if(rx_io_break) begin
      io_write_ready = 1'b1;
    end
  end

  assign io_write_thrown_payload = io_write_payload;
  assign io_write_thrown_ready = tx_io_write_ready;
  assign io_read_valid = rx_io_read_valid;
  assign io_read_payload = rx_io_read_payload;
  assign io_uart_txd = tx_io_txd;
  assign io_readError = rx_io_error;
  assign io_readBreak = rx_io_break;
  always @(posedge CLK_50 or posedge _zz_LED_R6) begin
    if(_zz_LED_R6) begin
      clockDivider_counter <= 20'h0;
      clockDivider_tickReg <= 1'b0;
    end else begin
      clockDivider_tickReg <= clockDivider_tick;
      clockDivider_counter <= (clockDivider_counter - 20'h00001);
      if(clockDivider_tick) begin
        clockDivider_counter <= io_config_clockDivider;
      end
    end
  end


endmodule

//UartCtrlRx_1 replaced by UartCtrlRx_1

//UartCtrlTx_1 replaced by UartCtrlTx_1

module Debounce (
  input      [102:0]  key_down,
  output              keyStatus_0_valid,
  output              keyStatus_0_payload,
  output              keyStatus_1_valid,
  output              keyStatus_1_payload,
  output              keyStatus_2_valid,
  output              keyStatus_2_payload,
  output              keyStatus_3_valid,
  output              keyStatus_3_payload,
  output              keyStatus_4_valid,
  output              keyStatus_4_payload,
  output              keyStatus_5_valid,
  output              keyStatus_5_payload,
  output              keyStatus_6_valid,
  output              keyStatus_6_payload,
  output              keyStatus_7_valid,
  output              keyStatus_7_payload,
  output              keyStatus_8_valid,
  output              keyStatus_8_payload,
  output              keyStatus_9_valid,
  output              keyStatus_9_payload,
  output              keyStatus_10_valid,
  output              keyStatus_10_payload,
  output              keyStatus_11_valid,
  output              keyStatus_11_payload,
  output              keyStatus_12_valid,
  output              keyStatus_12_payload,
  output              keyStatus_13_valid,
  output              keyStatus_13_payload,
  output              keyStatus_14_valid,
  output              keyStatus_14_payload,
  output              keyStatus_15_valid,
  output              keyStatus_15_payload,
  output              keyStatus_16_valid,
  output              keyStatus_16_payload,
  output              keyStatus_17_valid,
  output              keyStatus_17_payload,
  output              keyStatus_18_valid,
  output              keyStatus_18_payload,
  output              keyStatus_19_valid,
  output              keyStatus_19_payload,
  output              keyStatus_20_valid,
  output              keyStatus_20_payload,
  output              keyStatus_21_valid,
  output              keyStatus_21_payload,
  output              keyStatus_22_valid,
  output              keyStatus_22_payload,
  output              keyStatus_23_valid,
  output              keyStatus_23_payload,
  output              keyStatus_24_valid,
  output              keyStatus_24_payload,
  output              keyStatus_25_valid,
  output              keyStatus_25_payload,
  output              keyStatus_26_valid,
  output              keyStatus_26_payload,
  output              keyStatus_27_valid,
  output              keyStatus_27_payload,
  output              keyStatus_28_valid,
  output              keyStatus_28_payload,
  output              keyStatus_29_valid,
  output              keyStatus_29_payload,
  output              keyStatus_30_valid,
  output              keyStatus_30_payload,
  output              keyStatus_31_valid,
  output              keyStatus_31_payload,
  output              keyStatus_32_valid,
  output              keyStatus_32_payload,
  output              keyStatus_33_valid,
  output              keyStatus_33_payload,
  output              keyStatus_34_valid,
  output              keyStatus_34_payload,
  output              keyStatus_35_valid,
  output              keyStatus_35_payload,
  output              keyStatus_36_valid,
  output              keyStatus_36_payload,
  output              keyStatus_37_valid,
  output              keyStatus_37_payload,
  output              keyStatus_38_valid,
  output              keyStatus_38_payload,
  output              keyStatus_39_valid,
  output              keyStatus_39_payload,
  output              keyStatus_40_valid,
  output              keyStatus_40_payload,
  output              keyStatus_41_valid,
  output              keyStatus_41_payload,
  output              keyStatus_42_valid,
  output              keyStatus_42_payload,
  output              keyStatus_43_valid,
  output              keyStatus_43_payload,
  output              keyStatus_44_valid,
  output              keyStatus_44_payload,
  output              keyStatus_45_valid,
  output              keyStatus_45_payload,
  output              keyStatus_46_valid,
  output              keyStatus_46_payload,
  output              keyStatus_47_valid,
  output              keyStatus_47_payload,
  output              keyStatus_48_valid,
  output              keyStatus_48_payload,
  output              keyStatus_49_valid,
  output              keyStatus_49_payload,
  output              keyStatus_50_valid,
  output              keyStatus_50_payload,
  output              keyStatus_51_valid,
  output              keyStatus_51_payload,
  output              keyStatus_52_valid,
  output              keyStatus_52_payload,
  output              keyStatus_53_valid,
  output              keyStatus_53_payload,
  output              keyStatus_54_valid,
  output              keyStatus_54_payload,
  output              keyStatus_55_valid,
  output              keyStatus_55_payload,
  output              keyStatus_56_valid,
  output              keyStatus_56_payload,
  output              keyStatus_57_valid,
  output              keyStatus_57_payload,
  output              keyStatus_58_valid,
  output              keyStatus_58_payload,
  output              keyStatus_59_valid,
  output              keyStatus_59_payload,
  output              keyStatus_60_valid,
  output              keyStatus_60_payload,
  output              keyStatus_61_valid,
  output              keyStatus_61_payload,
  output              keyStatus_62_valid,
  output              keyStatus_62_payload,
  output              keyStatus_63_valid,
  output              keyStatus_63_payload,
  output              keyStatus_64_valid,
  output              keyStatus_64_payload,
  output              keyStatus_65_valid,
  output              keyStatus_65_payload,
  output              keyStatus_66_valid,
  output              keyStatus_66_payload,
  output              keyStatus_67_valid,
  output              keyStatus_67_payload,
  output              keyStatus_68_valid,
  output              keyStatus_68_payload,
  output              keyStatus_69_valid,
  output              keyStatus_69_payload,
  output              keyStatus_70_valid,
  output              keyStatus_70_payload,
  output              keyStatus_71_valid,
  output              keyStatus_71_payload,
  output              keyStatus_72_valid,
  output              keyStatus_72_payload,
  output              keyStatus_73_valid,
  output              keyStatus_73_payload,
  output              keyStatus_74_valid,
  output              keyStatus_74_payload,
  output              keyStatus_75_valid,
  output              keyStatus_75_payload,
  output              keyStatus_76_valid,
  output              keyStatus_76_payload,
  output              keyStatus_77_valid,
  output              keyStatus_77_payload,
  output              keyStatus_78_valid,
  output              keyStatus_78_payload,
  output              keyStatus_79_valid,
  output              keyStatus_79_payload,
  output              keyStatus_80_valid,
  output              keyStatus_80_payload,
  output              keyStatus_81_valid,
  output              keyStatus_81_payload,
  output              keyStatus_82_valid,
  output              keyStatus_82_payload,
  output              keyStatus_83_valid,
  output              keyStatus_83_payload,
  output              keyStatus_84_valid,
  output              keyStatus_84_payload,
  output              keyStatus_85_valid,
  output              keyStatus_85_payload,
  output              keyStatus_86_valid,
  output              keyStatus_86_payload,
  output              keyStatus_87_valid,
  output              keyStatus_87_payload,
  output              keyStatus_88_valid,
  output              keyStatus_88_payload,
  output              keyStatus_89_valid,
  output              keyStatus_89_payload,
  output              keyStatus_90_valid,
  output              keyStatus_90_payload,
  output              keyStatus_91_valid,
  output              keyStatus_91_payload,
  output              keyStatus_92_valid,
  output              keyStatus_92_payload,
  output              keyStatus_93_valid,
  output              keyStatus_93_payload,
  output              keyStatus_94_valid,
  output              keyStatus_94_payload,
  output              keyStatus_95_valid,
  output              keyStatus_95_payload,
  output              keyStatus_96_valid,
  output              keyStatus_96_payload,
  output              keyStatus_97_valid,
  output              keyStatus_97_payload,
  output              keyStatus_98_valid,
  output              keyStatus_98_payload,
  output              keyStatus_99_valid,
  output              keyStatus_99_payload,
  output              keyStatus_100_valid,
  output              keyStatus_100_payload,
  output              keyStatus_101_valid,
  output              keyStatus_101_payload,
  output              keyStatus_102_valid,
  output              keyStatus_102_payload,
  input               CLK_50,
  input               _zz_LED_R6
);

  wire                singleKey_103_raw;
  wire                singleKey_104_raw;
  wire                singleKey_105_raw;
  wire                singleKey_106_raw;
  wire                singleKey_107_raw;
  wire                singleKey_108_raw;
  wire                singleKey_109_raw;
  wire                singleKey_110_raw;
  wire                singleKey_111_raw;
  wire                singleKey_112_raw;
  wire                singleKey_113_raw;
  wire                singleKey_114_raw;
  wire                singleKey_115_raw;
  wire                singleKey_116_raw;
  wire                singleKey_117_raw;
  wire                singleKey_118_raw;
  wire                singleKey_119_raw;
  wire                singleKey_120_raw;
  wire                singleKey_121_raw;
  wire                singleKey_122_raw;
  wire                singleKey_123_raw;
  wire                singleKey_124_raw;
  wire                singleKey_125_raw;
  wire                singleKey_126_raw;
  wire                singleKey_127_raw;
  wire                singleKey_128_raw;
  wire                singleKey_129_raw;
  wire                singleKey_130_raw;
  wire                singleKey_131_raw;
  wire                singleKey_132_raw;
  wire                singleKey_133_raw;
  wire                singleKey_134_raw;
  wire                singleKey_135_raw;
  wire                singleKey_136_raw;
  wire                singleKey_137_raw;
  wire                singleKey_138_raw;
  wire                singleKey_139_raw;
  wire                singleKey_140_raw;
  wire                singleKey_141_raw;
  wire                singleKey_142_raw;
  wire                singleKey_143_raw;
  wire                singleKey_144_raw;
  wire                singleKey_145_raw;
  wire                singleKey_146_raw;
  wire                singleKey_147_raw;
  wire                singleKey_148_raw;
  wire                singleKey_149_raw;
  wire                singleKey_150_raw;
  wire                singleKey_151_raw;
  wire                singleKey_152_raw;
  wire                singleKey_153_raw;
  wire                singleKey_154_raw;
  wire                singleKey_155_raw;
  wire                singleKey_156_raw;
  wire                singleKey_157_raw;
  wire                singleKey_158_raw;
  wire                singleKey_159_raw;
  wire                singleKey_160_raw;
  wire                singleKey_161_raw;
  wire                singleKey_162_raw;
  wire                singleKey_163_raw;
  wire                singleKey_164_raw;
  wire                singleKey_165_raw;
  wire                singleKey_166_raw;
  wire                singleKey_167_raw;
  wire                singleKey_168_raw;
  wire                singleKey_169_raw;
  wire                singleKey_170_raw;
  wire                singleKey_171_raw;
  wire                singleKey_172_raw;
  wire                singleKey_173_raw;
  wire                singleKey_174_raw;
  wire                singleKey_175_raw;
  wire                singleKey_176_raw;
  wire                singleKey_177_raw;
  wire                singleKey_178_raw;
  wire                singleKey_179_raw;
  wire                singleKey_180_raw;
  wire                singleKey_181_raw;
  wire                singleKey_182_raw;
  wire                singleKey_183_raw;
  wire                singleKey_184_raw;
  wire                singleKey_185_raw;
  wire                singleKey_186_raw;
  wire                singleKey_187_raw;
  wire                singleKey_188_raw;
  wire                singleKey_189_raw;
  wire                singleKey_190_raw;
  wire                singleKey_191_raw;
  wire                singleKey_192_raw;
  wire                singleKey_193_raw;
  wire                singleKey_194_raw;
  wire                singleKey_195_raw;
  wire                singleKey_196_raw;
  wire                singleKey_197_raw;
  wire                singleKey_198_raw;
  wire                singleKey_199_raw;
  wire                singleKey_200_raw;
  wire                singleKey_201_raw;
  wire                singleKey_202_raw;
  wire                singleKey_203_raw;
  wire                singleKey_204_raw;
  wire                singleKey_205_raw;
  wire                singleKey_103_filtered_valid;
  wire                singleKey_103_filtered_payload;
  wire                singleKey_104_filtered_valid;
  wire                singleKey_104_filtered_payload;
  wire                singleKey_105_filtered_valid;
  wire                singleKey_105_filtered_payload;
  wire                singleKey_106_filtered_valid;
  wire                singleKey_106_filtered_payload;
  wire                singleKey_107_filtered_valid;
  wire                singleKey_107_filtered_payload;
  wire                singleKey_108_filtered_valid;
  wire                singleKey_108_filtered_payload;
  wire                singleKey_109_filtered_valid;
  wire                singleKey_109_filtered_payload;
  wire                singleKey_110_filtered_valid;
  wire                singleKey_110_filtered_payload;
  wire                singleKey_111_filtered_valid;
  wire                singleKey_111_filtered_payload;
  wire                singleKey_112_filtered_valid;
  wire                singleKey_112_filtered_payload;
  wire                singleKey_113_filtered_valid;
  wire                singleKey_113_filtered_payload;
  wire                singleKey_114_filtered_valid;
  wire                singleKey_114_filtered_payload;
  wire                singleKey_115_filtered_valid;
  wire                singleKey_115_filtered_payload;
  wire                singleKey_116_filtered_valid;
  wire                singleKey_116_filtered_payload;
  wire                singleKey_117_filtered_valid;
  wire                singleKey_117_filtered_payload;
  wire                singleKey_118_filtered_valid;
  wire                singleKey_118_filtered_payload;
  wire                singleKey_119_filtered_valid;
  wire                singleKey_119_filtered_payload;
  wire                singleKey_120_filtered_valid;
  wire                singleKey_120_filtered_payload;
  wire                singleKey_121_filtered_valid;
  wire                singleKey_121_filtered_payload;
  wire                singleKey_122_filtered_valid;
  wire                singleKey_122_filtered_payload;
  wire                singleKey_123_filtered_valid;
  wire                singleKey_123_filtered_payload;
  wire                singleKey_124_filtered_valid;
  wire                singleKey_124_filtered_payload;
  wire                singleKey_125_filtered_valid;
  wire                singleKey_125_filtered_payload;
  wire                singleKey_126_filtered_valid;
  wire                singleKey_126_filtered_payload;
  wire                singleKey_127_filtered_valid;
  wire                singleKey_127_filtered_payload;
  wire                singleKey_128_filtered_valid;
  wire                singleKey_128_filtered_payload;
  wire                singleKey_129_filtered_valid;
  wire                singleKey_129_filtered_payload;
  wire                singleKey_130_filtered_valid;
  wire                singleKey_130_filtered_payload;
  wire                singleKey_131_filtered_valid;
  wire                singleKey_131_filtered_payload;
  wire                singleKey_132_filtered_valid;
  wire                singleKey_132_filtered_payload;
  wire                singleKey_133_filtered_valid;
  wire                singleKey_133_filtered_payload;
  wire                singleKey_134_filtered_valid;
  wire                singleKey_134_filtered_payload;
  wire                singleKey_135_filtered_valid;
  wire                singleKey_135_filtered_payload;
  wire                singleKey_136_filtered_valid;
  wire                singleKey_136_filtered_payload;
  wire                singleKey_137_filtered_valid;
  wire                singleKey_137_filtered_payload;
  wire                singleKey_138_filtered_valid;
  wire                singleKey_138_filtered_payload;
  wire                singleKey_139_filtered_valid;
  wire                singleKey_139_filtered_payload;
  wire                singleKey_140_filtered_valid;
  wire                singleKey_140_filtered_payload;
  wire                singleKey_141_filtered_valid;
  wire                singleKey_141_filtered_payload;
  wire                singleKey_142_filtered_valid;
  wire                singleKey_142_filtered_payload;
  wire                singleKey_143_filtered_valid;
  wire                singleKey_143_filtered_payload;
  wire                singleKey_144_filtered_valid;
  wire                singleKey_144_filtered_payload;
  wire                singleKey_145_filtered_valid;
  wire                singleKey_145_filtered_payload;
  wire                singleKey_146_filtered_valid;
  wire                singleKey_146_filtered_payload;
  wire                singleKey_147_filtered_valid;
  wire                singleKey_147_filtered_payload;
  wire                singleKey_148_filtered_valid;
  wire                singleKey_148_filtered_payload;
  wire                singleKey_149_filtered_valid;
  wire                singleKey_149_filtered_payload;
  wire                singleKey_150_filtered_valid;
  wire                singleKey_150_filtered_payload;
  wire                singleKey_151_filtered_valid;
  wire                singleKey_151_filtered_payload;
  wire                singleKey_152_filtered_valid;
  wire                singleKey_152_filtered_payload;
  wire                singleKey_153_filtered_valid;
  wire                singleKey_153_filtered_payload;
  wire                singleKey_154_filtered_valid;
  wire                singleKey_154_filtered_payload;
  wire                singleKey_155_filtered_valid;
  wire                singleKey_155_filtered_payload;
  wire                singleKey_156_filtered_valid;
  wire                singleKey_156_filtered_payload;
  wire                singleKey_157_filtered_valid;
  wire                singleKey_157_filtered_payload;
  wire                singleKey_158_filtered_valid;
  wire                singleKey_158_filtered_payload;
  wire                singleKey_159_filtered_valid;
  wire                singleKey_159_filtered_payload;
  wire                singleKey_160_filtered_valid;
  wire                singleKey_160_filtered_payload;
  wire                singleKey_161_filtered_valid;
  wire                singleKey_161_filtered_payload;
  wire                singleKey_162_filtered_valid;
  wire                singleKey_162_filtered_payload;
  wire                singleKey_163_filtered_valid;
  wire                singleKey_163_filtered_payload;
  wire                singleKey_164_filtered_valid;
  wire                singleKey_164_filtered_payload;
  wire                singleKey_165_filtered_valid;
  wire                singleKey_165_filtered_payload;
  wire                singleKey_166_filtered_valid;
  wire                singleKey_166_filtered_payload;
  wire                singleKey_167_filtered_valid;
  wire                singleKey_167_filtered_payload;
  wire                singleKey_168_filtered_valid;
  wire                singleKey_168_filtered_payload;
  wire                singleKey_169_filtered_valid;
  wire                singleKey_169_filtered_payload;
  wire                singleKey_170_filtered_valid;
  wire                singleKey_170_filtered_payload;
  wire                singleKey_171_filtered_valid;
  wire                singleKey_171_filtered_payload;
  wire                singleKey_172_filtered_valid;
  wire                singleKey_172_filtered_payload;
  wire                singleKey_173_filtered_valid;
  wire                singleKey_173_filtered_payload;
  wire                singleKey_174_filtered_valid;
  wire                singleKey_174_filtered_payload;
  wire                singleKey_175_filtered_valid;
  wire                singleKey_175_filtered_payload;
  wire                singleKey_176_filtered_valid;
  wire                singleKey_176_filtered_payload;
  wire                singleKey_177_filtered_valid;
  wire                singleKey_177_filtered_payload;
  wire                singleKey_178_filtered_valid;
  wire                singleKey_178_filtered_payload;
  wire                singleKey_179_filtered_valid;
  wire                singleKey_179_filtered_payload;
  wire                singleKey_180_filtered_valid;
  wire                singleKey_180_filtered_payload;
  wire                singleKey_181_filtered_valid;
  wire                singleKey_181_filtered_payload;
  wire                singleKey_182_filtered_valid;
  wire                singleKey_182_filtered_payload;
  wire                singleKey_183_filtered_valid;
  wire                singleKey_183_filtered_payload;
  wire                singleKey_184_filtered_valid;
  wire                singleKey_184_filtered_payload;
  wire                singleKey_185_filtered_valid;
  wire                singleKey_185_filtered_payload;
  wire                singleKey_186_filtered_valid;
  wire                singleKey_186_filtered_payload;
  wire                singleKey_187_filtered_valid;
  wire                singleKey_187_filtered_payload;
  wire                singleKey_188_filtered_valid;
  wire                singleKey_188_filtered_payload;
  wire                singleKey_189_filtered_valid;
  wire                singleKey_189_filtered_payload;
  wire                singleKey_190_filtered_valid;
  wire                singleKey_190_filtered_payload;
  wire                singleKey_191_filtered_valid;
  wire                singleKey_191_filtered_payload;
  wire                singleKey_192_filtered_valid;
  wire                singleKey_192_filtered_payload;
  wire                singleKey_193_filtered_valid;
  wire                singleKey_193_filtered_payload;
  wire                singleKey_194_filtered_valid;
  wire                singleKey_194_filtered_payload;
  wire                singleKey_195_filtered_valid;
  wire                singleKey_195_filtered_payload;
  wire                singleKey_196_filtered_valid;
  wire                singleKey_196_filtered_payload;
  wire                singleKey_197_filtered_valid;
  wire                singleKey_197_filtered_payload;
  wire                singleKey_198_filtered_valid;
  wire                singleKey_198_filtered_payload;
  wire                singleKey_199_filtered_valid;
  wire                singleKey_199_filtered_payload;
  wire                singleKey_200_filtered_valid;
  wire                singleKey_200_filtered_payload;
  wire                singleKey_201_filtered_valid;
  wire                singleKey_201_filtered_payload;
  wire                singleKey_202_filtered_valid;
  wire                singleKey_202_filtered_payload;
  wire                singleKey_203_filtered_valid;
  wire                singleKey_203_filtered_payload;
  wire                singleKey_204_filtered_valid;
  wire                singleKey_204_filtered_payload;
  wire                singleKey_205_filtered_valid;
  wire                singleKey_205_filtered_payload;
  reg        [14:0]   _zz_when_ClockDomain_l369;
  wire                when_ClockDomain_l369;
  reg                 when_ClockDomain_l369_regNext;

  SingleKey_102 singleKey_103 (
    .raw                           (singleKey_103_raw             ), //i
    .filtered_valid                (singleKey_103_filtered_valid  ), //o
    .filtered_payload              (singleKey_103_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_104 (
    .raw                           (singleKey_104_raw             ), //i
    .filtered_valid                (singleKey_104_filtered_valid  ), //o
    .filtered_payload              (singleKey_104_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_105 (
    .raw                           (singleKey_105_raw             ), //i
    .filtered_valid                (singleKey_105_filtered_valid  ), //o
    .filtered_payload              (singleKey_105_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_106 (
    .raw                           (singleKey_106_raw             ), //i
    .filtered_valid                (singleKey_106_filtered_valid  ), //o
    .filtered_payload              (singleKey_106_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_107 (
    .raw                           (singleKey_107_raw             ), //i
    .filtered_valid                (singleKey_107_filtered_valid  ), //o
    .filtered_payload              (singleKey_107_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_108 (
    .raw                           (singleKey_108_raw             ), //i
    .filtered_valid                (singleKey_108_filtered_valid  ), //o
    .filtered_payload              (singleKey_108_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_109 (
    .raw                           (singleKey_109_raw             ), //i
    .filtered_valid                (singleKey_109_filtered_valid  ), //o
    .filtered_payload              (singleKey_109_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_110 (
    .raw                           (singleKey_110_raw             ), //i
    .filtered_valid                (singleKey_110_filtered_valid  ), //o
    .filtered_payload              (singleKey_110_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_111 (
    .raw                           (singleKey_111_raw             ), //i
    .filtered_valid                (singleKey_111_filtered_valid  ), //o
    .filtered_payload              (singleKey_111_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_112 (
    .raw                           (singleKey_112_raw             ), //i
    .filtered_valid                (singleKey_112_filtered_valid  ), //o
    .filtered_payload              (singleKey_112_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_113 (
    .raw                           (singleKey_113_raw             ), //i
    .filtered_valid                (singleKey_113_filtered_valid  ), //o
    .filtered_payload              (singleKey_113_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_114 (
    .raw                           (singleKey_114_raw             ), //i
    .filtered_valid                (singleKey_114_filtered_valid  ), //o
    .filtered_payload              (singleKey_114_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_115 (
    .raw                           (singleKey_115_raw             ), //i
    .filtered_valid                (singleKey_115_filtered_valid  ), //o
    .filtered_payload              (singleKey_115_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_116 (
    .raw                           (singleKey_116_raw             ), //i
    .filtered_valid                (singleKey_116_filtered_valid  ), //o
    .filtered_payload              (singleKey_116_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_117 (
    .raw                           (singleKey_117_raw             ), //i
    .filtered_valid                (singleKey_117_filtered_valid  ), //o
    .filtered_payload              (singleKey_117_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_118 (
    .raw                           (singleKey_118_raw             ), //i
    .filtered_valid                (singleKey_118_filtered_valid  ), //o
    .filtered_payload              (singleKey_118_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_119 (
    .raw                           (singleKey_119_raw             ), //i
    .filtered_valid                (singleKey_119_filtered_valid  ), //o
    .filtered_payload              (singleKey_119_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_120 (
    .raw                           (singleKey_120_raw             ), //i
    .filtered_valid                (singleKey_120_filtered_valid  ), //o
    .filtered_payload              (singleKey_120_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_121 (
    .raw                           (singleKey_121_raw             ), //i
    .filtered_valid                (singleKey_121_filtered_valid  ), //o
    .filtered_payload              (singleKey_121_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_122 (
    .raw                           (singleKey_122_raw             ), //i
    .filtered_valid                (singleKey_122_filtered_valid  ), //o
    .filtered_payload              (singleKey_122_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_123 (
    .raw                           (singleKey_123_raw             ), //i
    .filtered_valid                (singleKey_123_filtered_valid  ), //o
    .filtered_payload              (singleKey_123_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_124 (
    .raw                           (singleKey_124_raw             ), //i
    .filtered_valid                (singleKey_124_filtered_valid  ), //o
    .filtered_payload              (singleKey_124_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_125 (
    .raw                           (singleKey_125_raw             ), //i
    .filtered_valid                (singleKey_125_filtered_valid  ), //o
    .filtered_payload              (singleKey_125_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_126 (
    .raw                           (singleKey_126_raw             ), //i
    .filtered_valid                (singleKey_126_filtered_valid  ), //o
    .filtered_payload              (singleKey_126_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_127 (
    .raw                           (singleKey_127_raw             ), //i
    .filtered_valid                (singleKey_127_filtered_valid  ), //o
    .filtered_payload              (singleKey_127_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_128 (
    .raw                           (singleKey_128_raw             ), //i
    .filtered_valid                (singleKey_128_filtered_valid  ), //o
    .filtered_payload              (singleKey_128_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_129 (
    .raw                           (singleKey_129_raw             ), //i
    .filtered_valid                (singleKey_129_filtered_valid  ), //o
    .filtered_payload              (singleKey_129_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_130 (
    .raw                           (singleKey_130_raw             ), //i
    .filtered_valid                (singleKey_130_filtered_valid  ), //o
    .filtered_payload              (singleKey_130_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_131 (
    .raw                           (singleKey_131_raw             ), //i
    .filtered_valid                (singleKey_131_filtered_valid  ), //o
    .filtered_payload              (singleKey_131_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_132 (
    .raw                           (singleKey_132_raw             ), //i
    .filtered_valid                (singleKey_132_filtered_valid  ), //o
    .filtered_payload              (singleKey_132_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_133 (
    .raw                           (singleKey_133_raw             ), //i
    .filtered_valid                (singleKey_133_filtered_valid  ), //o
    .filtered_payload              (singleKey_133_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_134 (
    .raw                           (singleKey_134_raw             ), //i
    .filtered_valid                (singleKey_134_filtered_valid  ), //o
    .filtered_payload              (singleKey_134_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_135 (
    .raw                           (singleKey_135_raw             ), //i
    .filtered_valid                (singleKey_135_filtered_valid  ), //o
    .filtered_payload              (singleKey_135_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_136 (
    .raw                           (singleKey_136_raw             ), //i
    .filtered_valid                (singleKey_136_filtered_valid  ), //o
    .filtered_payload              (singleKey_136_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_137 (
    .raw                           (singleKey_137_raw             ), //i
    .filtered_valid                (singleKey_137_filtered_valid  ), //o
    .filtered_payload              (singleKey_137_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_138 (
    .raw                           (singleKey_138_raw             ), //i
    .filtered_valid                (singleKey_138_filtered_valid  ), //o
    .filtered_payload              (singleKey_138_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_139 (
    .raw                           (singleKey_139_raw             ), //i
    .filtered_valid                (singleKey_139_filtered_valid  ), //o
    .filtered_payload              (singleKey_139_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_140 (
    .raw                           (singleKey_140_raw             ), //i
    .filtered_valid                (singleKey_140_filtered_valid  ), //o
    .filtered_payload              (singleKey_140_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_141 (
    .raw                           (singleKey_141_raw             ), //i
    .filtered_valid                (singleKey_141_filtered_valid  ), //o
    .filtered_payload              (singleKey_141_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_142 (
    .raw                           (singleKey_142_raw             ), //i
    .filtered_valid                (singleKey_142_filtered_valid  ), //o
    .filtered_payload              (singleKey_142_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_143 (
    .raw                           (singleKey_143_raw             ), //i
    .filtered_valid                (singleKey_143_filtered_valid  ), //o
    .filtered_payload              (singleKey_143_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_144 (
    .raw                           (singleKey_144_raw             ), //i
    .filtered_valid                (singleKey_144_filtered_valid  ), //o
    .filtered_payload              (singleKey_144_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_145 (
    .raw                           (singleKey_145_raw             ), //i
    .filtered_valid                (singleKey_145_filtered_valid  ), //o
    .filtered_payload              (singleKey_145_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_146 (
    .raw                           (singleKey_146_raw             ), //i
    .filtered_valid                (singleKey_146_filtered_valid  ), //o
    .filtered_payload              (singleKey_146_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_147 (
    .raw                           (singleKey_147_raw             ), //i
    .filtered_valid                (singleKey_147_filtered_valid  ), //o
    .filtered_payload              (singleKey_147_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_148 (
    .raw                           (singleKey_148_raw             ), //i
    .filtered_valid                (singleKey_148_filtered_valid  ), //o
    .filtered_payload              (singleKey_148_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_149 (
    .raw                           (singleKey_149_raw             ), //i
    .filtered_valid                (singleKey_149_filtered_valid  ), //o
    .filtered_payload              (singleKey_149_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_150 (
    .raw                           (singleKey_150_raw             ), //i
    .filtered_valid                (singleKey_150_filtered_valid  ), //o
    .filtered_payload              (singleKey_150_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_151 (
    .raw                           (singleKey_151_raw             ), //i
    .filtered_valid                (singleKey_151_filtered_valid  ), //o
    .filtered_payload              (singleKey_151_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_152 (
    .raw                           (singleKey_152_raw             ), //i
    .filtered_valid                (singleKey_152_filtered_valid  ), //o
    .filtered_payload              (singleKey_152_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_153 (
    .raw                           (singleKey_153_raw             ), //i
    .filtered_valid                (singleKey_153_filtered_valid  ), //o
    .filtered_payload              (singleKey_153_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_154 (
    .raw                           (singleKey_154_raw             ), //i
    .filtered_valid                (singleKey_154_filtered_valid  ), //o
    .filtered_payload              (singleKey_154_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_155 (
    .raw                           (singleKey_155_raw             ), //i
    .filtered_valid                (singleKey_155_filtered_valid  ), //o
    .filtered_payload              (singleKey_155_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_156 (
    .raw                           (singleKey_156_raw             ), //i
    .filtered_valid                (singleKey_156_filtered_valid  ), //o
    .filtered_payload              (singleKey_156_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_157 (
    .raw                           (singleKey_157_raw             ), //i
    .filtered_valid                (singleKey_157_filtered_valid  ), //o
    .filtered_payload              (singleKey_157_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_158 (
    .raw                           (singleKey_158_raw             ), //i
    .filtered_valid                (singleKey_158_filtered_valid  ), //o
    .filtered_payload              (singleKey_158_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_159 (
    .raw                           (singleKey_159_raw             ), //i
    .filtered_valid                (singleKey_159_filtered_valid  ), //o
    .filtered_payload              (singleKey_159_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_160 (
    .raw                           (singleKey_160_raw             ), //i
    .filtered_valid                (singleKey_160_filtered_valid  ), //o
    .filtered_payload              (singleKey_160_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_161 (
    .raw                           (singleKey_161_raw             ), //i
    .filtered_valid                (singleKey_161_filtered_valid  ), //o
    .filtered_payload              (singleKey_161_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_162 (
    .raw                           (singleKey_162_raw             ), //i
    .filtered_valid                (singleKey_162_filtered_valid  ), //o
    .filtered_payload              (singleKey_162_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_163 (
    .raw                           (singleKey_163_raw             ), //i
    .filtered_valid                (singleKey_163_filtered_valid  ), //o
    .filtered_payload              (singleKey_163_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_164 (
    .raw                           (singleKey_164_raw             ), //i
    .filtered_valid                (singleKey_164_filtered_valid  ), //o
    .filtered_payload              (singleKey_164_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_165 (
    .raw                           (singleKey_165_raw             ), //i
    .filtered_valid                (singleKey_165_filtered_valid  ), //o
    .filtered_payload              (singleKey_165_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_166 (
    .raw                           (singleKey_166_raw             ), //i
    .filtered_valid                (singleKey_166_filtered_valid  ), //o
    .filtered_payload              (singleKey_166_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_167 (
    .raw                           (singleKey_167_raw             ), //i
    .filtered_valid                (singleKey_167_filtered_valid  ), //o
    .filtered_payload              (singleKey_167_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_168 (
    .raw                           (singleKey_168_raw             ), //i
    .filtered_valid                (singleKey_168_filtered_valid  ), //o
    .filtered_payload              (singleKey_168_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_169 (
    .raw                           (singleKey_169_raw             ), //i
    .filtered_valid                (singleKey_169_filtered_valid  ), //o
    .filtered_payload              (singleKey_169_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_170 (
    .raw                           (singleKey_170_raw             ), //i
    .filtered_valid                (singleKey_170_filtered_valid  ), //o
    .filtered_payload              (singleKey_170_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_171 (
    .raw                           (singleKey_171_raw             ), //i
    .filtered_valid                (singleKey_171_filtered_valid  ), //o
    .filtered_payload              (singleKey_171_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_172 (
    .raw                           (singleKey_172_raw             ), //i
    .filtered_valid                (singleKey_172_filtered_valid  ), //o
    .filtered_payload              (singleKey_172_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_173 (
    .raw                           (singleKey_173_raw             ), //i
    .filtered_valid                (singleKey_173_filtered_valid  ), //o
    .filtered_payload              (singleKey_173_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_174 (
    .raw                           (singleKey_174_raw             ), //i
    .filtered_valid                (singleKey_174_filtered_valid  ), //o
    .filtered_payload              (singleKey_174_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_175 (
    .raw                           (singleKey_175_raw             ), //i
    .filtered_valid                (singleKey_175_filtered_valid  ), //o
    .filtered_payload              (singleKey_175_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_176 (
    .raw                           (singleKey_176_raw             ), //i
    .filtered_valid                (singleKey_176_filtered_valid  ), //o
    .filtered_payload              (singleKey_176_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_177 (
    .raw                           (singleKey_177_raw             ), //i
    .filtered_valid                (singleKey_177_filtered_valid  ), //o
    .filtered_payload              (singleKey_177_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_178 (
    .raw                           (singleKey_178_raw             ), //i
    .filtered_valid                (singleKey_178_filtered_valid  ), //o
    .filtered_payload              (singleKey_178_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_179 (
    .raw                           (singleKey_179_raw             ), //i
    .filtered_valid                (singleKey_179_filtered_valid  ), //o
    .filtered_payload              (singleKey_179_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_180 (
    .raw                           (singleKey_180_raw             ), //i
    .filtered_valid                (singleKey_180_filtered_valid  ), //o
    .filtered_payload              (singleKey_180_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_181 (
    .raw                           (singleKey_181_raw             ), //i
    .filtered_valid                (singleKey_181_filtered_valid  ), //o
    .filtered_payload              (singleKey_181_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_182 (
    .raw                           (singleKey_182_raw             ), //i
    .filtered_valid                (singleKey_182_filtered_valid  ), //o
    .filtered_payload              (singleKey_182_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_183 (
    .raw                           (singleKey_183_raw             ), //i
    .filtered_valid                (singleKey_183_filtered_valid  ), //o
    .filtered_payload              (singleKey_183_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_184 (
    .raw                           (singleKey_184_raw             ), //i
    .filtered_valid                (singleKey_184_filtered_valid  ), //o
    .filtered_payload              (singleKey_184_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_185 (
    .raw                           (singleKey_185_raw             ), //i
    .filtered_valid                (singleKey_185_filtered_valid  ), //o
    .filtered_payload              (singleKey_185_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_186 (
    .raw                           (singleKey_186_raw             ), //i
    .filtered_valid                (singleKey_186_filtered_valid  ), //o
    .filtered_payload              (singleKey_186_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_187 (
    .raw                           (singleKey_187_raw             ), //i
    .filtered_valid                (singleKey_187_filtered_valid  ), //o
    .filtered_payload              (singleKey_187_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_188 (
    .raw                           (singleKey_188_raw             ), //i
    .filtered_valid                (singleKey_188_filtered_valid  ), //o
    .filtered_payload              (singleKey_188_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_189 (
    .raw                           (singleKey_189_raw             ), //i
    .filtered_valid                (singleKey_189_filtered_valid  ), //o
    .filtered_payload              (singleKey_189_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_190 (
    .raw                           (singleKey_190_raw             ), //i
    .filtered_valid                (singleKey_190_filtered_valid  ), //o
    .filtered_payload              (singleKey_190_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_191 (
    .raw                           (singleKey_191_raw             ), //i
    .filtered_valid                (singleKey_191_filtered_valid  ), //o
    .filtered_payload              (singleKey_191_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_192 (
    .raw                           (singleKey_192_raw             ), //i
    .filtered_valid                (singleKey_192_filtered_valid  ), //o
    .filtered_payload              (singleKey_192_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_193 (
    .raw                           (singleKey_193_raw             ), //i
    .filtered_valid                (singleKey_193_filtered_valid  ), //o
    .filtered_payload              (singleKey_193_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_194 (
    .raw                           (singleKey_194_raw             ), //i
    .filtered_valid                (singleKey_194_filtered_valid  ), //o
    .filtered_payload              (singleKey_194_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_195 (
    .raw                           (singleKey_195_raw             ), //i
    .filtered_valid                (singleKey_195_filtered_valid  ), //o
    .filtered_payload              (singleKey_195_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_196 (
    .raw                           (singleKey_196_raw             ), //i
    .filtered_valid                (singleKey_196_filtered_valid  ), //o
    .filtered_payload              (singleKey_196_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_197 (
    .raw                           (singleKey_197_raw             ), //i
    .filtered_valid                (singleKey_197_filtered_valid  ), //o
    .filtered_payload              (singleKey_197_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_198 (
    .raw                           (singleKey_198_raw             ), //i
    .filtered_valid                (singleKey_198_filtered_valid  ), //o
    .filtered_payload              (singleKey_198_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_199 (
    .raw                           (singleKey_199_raw             ), //i
    .filtered_valid                (singleKey_199_filtered_valid  ), //o
    .filtered_payload              (singleKey_199_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_200 (
    .raw                           (singleKey_200_raw             ), //i
    .filtered_valid                (singleKey_200_filtered_valid  ), //o
    .filtered_payload              (singleKey_200_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_201 (
    .raw                           (singleKey_201_raw             ), //i
    .filtered_valid                (singleKey_201_filtered_valid  ), //o
    .filtered_payload              (singleKey_201_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_202 (
    .raw                           (singleKey_202_raw             ), //i
    .filtered_valid                (singleKey_202_filtered_valid  ), //o
    .filtered_payload              (singleKey_202_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_203 (
    .raw                           (singleKey_203_raw             ), //i
    .filtered_valid                (singleKey_203_filtered_valid  ), //o
    .filtered_payload              (singleKey_203_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_204 (
    .raw                           (singleKey_204_raw             ), //i
    .filtered_valid                (singleKey_204_filtered_valid  ), //o
    .filtered_payload              (singleKey_204_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  SingleKey_102 singleKey_205 (
    .raw                           (singleKey_205_raw             ), //i
    .filtered_valid                (singleKey_205_filtered_valid  ), //o
    .filtered_payload              (singleKey_205_filtered_payload), //o
    .CLK_50                        (CLK_50                        ), //i
    ._zz_LED_R6                    (_zz_LED_R6                    ), //i
    .when_ClockDomain_l369_regNext (when_ClockDomain_l369_regNext )  //i
  );
  assign when_ClockDomain_l369 = (_zz_when_ClockDomain_l369 == 15'h61a7);
  assign singleKey_103_raw = key_down[0];
  assign keyStatus_0_valid = singleKey_103_filtered_valid;
  assign keyStatus_0_payload = singleKey_103_filtered_payload;
  assign singleKey_104_raw = key_down[1];
  assign keyStatus_1_valid = singleKey_104_filtered_valid;
  assign keyStatus_1_payload = singleKey_104_filtered_payload;
  assign singleKey_105_raw = key_down[2];
  assign keyStatus_2_valid = singleKey_105_filtered_valid;
  assign keyStatus_2_payload = singleKey_105_filtered_payload;
  assign singleKey_106_raw = key_down[3];
  assign keyStatus_3_valid = singleKey_106_filtered_valid;
  assign keyStatus_3_payload = singleKey_106_filtered_payload;
  assign singleKey_107_raw = key_down[4];
  assign keyStatus_4_valid = singleKey_107_filtered_valid;
  assign keyStatus_4_payload = singleKey_107_filtered_payload;
  assign singleKey_108_raw = key_down[5];
  assign keyStatus_5_valid = singleKey_108_filtered_valid;
  assign keyStatus_5_payload = singleKey_108_filtered_payload;
  assign singleKey_109_raw = key_down[6];
  assign keyStatus_6_valid = singleKey_109_filtered_valid;
  assign keyStatus_6_payload = singleKey_109_filtered_payload;
  assign singleKey_110_raw = key_down[7];
  assign keyStatus_7_valid = singleKey_110_filtered_valid;
  assign keyStatus_7_payload = singleKey_110_filtered_payload;
  assign singleKey_111_raw = key_down[8];
  assign keyStatus_8_valid = singleKey_111_filtered_valid;
  assign keyStatus_8_payload = singleKey_111_filtered_payload;
  assign singleKey_112_raw = key_down[9];
  assign keyStatus_9_valid = singleKey_112_filtered_valid;
  assign keyStatus_9_payload = singleKey_112_filtered_payload;
  assign singleKey_113_raw = key_down[10];
  assign keyStatus_10_valid = singleKey_113_filtered_valid;
  assign keyStatus_10_payload = singleKey_113_filtered_payload;
  assign singleKey_114_raw = key_down[11];
  assign keyStatus_11_valid = singleKey_114_filtered_valid;
  assign keyStatus_11_payload = singleKey_114_filtered_payload;
  assign singleKey_115_raw = key_down[12];
  assign keyStatus_12_valid = singleKey_115_filtered_valid;
  assign keyStatus_12_payload = singleKey_115_filtered_payload;
  assign singleKey_116_raw = key_down[13];
  assign keyStatus_13_valid = singleKey_116_filtered_valid;
  assign keyStatus_13_payload = singleKey_116_filtered_payload;
  assign singleKey_117_raw = key_down[14];
  assign keyStatus_14_valid = singleKey_117_filtered_valid;
  assign keyStatus_14_payload = singleKey_117_filtered_payload;
  assign singleKey_118_raw = key_down[15];
  assign keyStatus_15_valid = singleKey_118_filtered_valid;
  assign keyStatus_15_payload = singleKey_118_filtered_payload;
  assign singleKey_119_raw = key_down[16];
  assign keyStatus_16_valid = singleKey_119_filtered_valid;
  assign keyStatus_16_payload = singleKey_119_filtered_payload;
  assign singleKey_120_raw = key_down[17];
  assign keyStatus_17_valid = singleKey_120_filtered_valid;
  assign keyStatus_17_payload = singleKey_120_filtered_payload;
  assign singleKey_121_raw = key_down[18];
  assign keyStatus_18_valid = singleKey_121_filtered_valid;
  assign keyStatus_18_payload = singleKey_121_filtered_payload;
  assign singleKey_122_raw = key_down[19];
  assign keyStatus_19_valid = singleKey_122_filtered_valid;
  assign keyStatus_19_payload = singleKey_122_filtered_payload;
  assign singleKey_123_raw = key_down[20];
  assign keyStatus_20_valid = singleKey_123_filtered_valid;
  assign keyStatus_20_payload = singleKey_123_filtered_payload;
  assign singleKey_124_raw = key_down[21];
  assign keyStatus_21_valid = singleKey_124_filtered_valid;
  assign keyStatus_21_payload = singleKey_124_filtered_payload;
  assign singleKey_125_raw = key_down[22];
  assign keyStatus_22_valid = singleKey_125_filtered_valid;
  assign keyStatus_22_payload = singleKey_125_filtered_payload;
  assign singleKey_126_raw = key_down[23];
  assign keyStatus_23_valid = singleKey_126_filtered_valid;
  assign keyStatus_23_payload = singleKey_126_filtered_payload;
  assign singleKey_127_raw = key_down[24];
  assign keyStatus_24_valid = singleKey_127_filtered_valid;
  assign keyStatus_24_payload = singleKey_127_filtered_payload;
  assign singleKey_128_raw = key_down[25];
  assign keyStatus_25_valid = singleKey_128_filtered_valid;
  assign keyStatus_25_payload = singleKey_128_filtered_payload;
  assign singleKey_129_raw = key_down[26];
  assign keyStatus_26_valid = singleKey_129_filtered_valid;
  assign keyStatus_26_payload = singleKey_129_filtered_payload;
  assign singleKey_130_raw = key_down[27];
  assign keyStatus_27_valid = singleKey_130_filtered_valid;
  assign keyStatus_27_payload = singleKey_130_filtered_payload;
  assign singleKey_131_raw = key_down[28];
  assign keyStatus_28_valid = singleKey_131_filtered_valid;
  assign keyStatus_28_payload = singleKey_131_filtered_payload;
  assign singleKey_132_raw = key_down[29];
  assign keyStatus_29_valid = singleKey_132_filtered_valid;
  assign keyStatus_29_payload = singleKey_132_filtered_payload;
  assign singleKey_133_raw = key_down[30];
  assign keyStatus_30_valid = singleKey_133_filtered_valid;
  assign keyStatus_30_payload = singleKey_133_filtered_payload;
  assign singleKey_134_raw = key_down[31];
  assign keyStatus_31_valid = singleKey_134_filtered_valid;
  assign keyStatus_31_payload = singleKey_134_filtered_payload;
  assign singleKey_135_raw = key_down[32];
  assign keyStatus_32_valid = singleKey_135_filtered_valid;
  assign keyStatus_32_payload = singleKey_135_filtered_payload;
  assign singleKey_136_raw = key_down[33];
  assign keyStatus_33_valid = singleKey_136_filtered_valid;
  assign keyStatus_33_payload = singleKey_136_filtered_payload;
  assign singleKey_137_raw = key_down[34];
  assign keyStatus_34_valid = singleKey_137_filtered_valid;
  assign keyStatus_34_payload = singleKey_137_filtered_payload;
  assign singleKey_138_raw = key_down[35];
  assign keyStatus_35_valid = singleKey_138_filtered_valid;
  assign keyStatus_35_payload = singleKey_138_filtered_payload;
  assign singleKey_139_raw = key_down[36];
  assign keyStatus_36_valid = singleKey_139_filtered_valid;
  assign keyStatus_36_payload = singleKey_139_filtered_payload;
  assign singleKey_140_raw = key_down[37];
  assign keyStatus_37_valid = singleKey_140_filtered_valid;
  assign keyStatus_37_payload = singleKey_140_filtered_payload;
  assign singleKey_141_raw = key_down[38];
  assign keyStatus_38_valid = singleKey_141_filtered_valid;
  assign keyStatus_38_payload = singleKey_141_filtered_payload;
  assign singleKey_142_raw = key_down[39];
  assign keyStatus_39_valid = singleKey_142_filtered_valid;
  assign keyStatus_39_payload = singleKey_142_filtered_payload;
  assign singleKey_143_raw = key_down[40];
  assign keyStatus_40_valid = singleKey_143_filtered_valid;
  assign keyStatus_40_payload = singleKey_143_filtered_payload;
  assign singleKey_144_raw = key_down[41];
  assign keyStatus_41_valid = singleKey_144_filtered_valid;
  assign keyStatus_41_payload = singleKey_144_filtered_payload;
  assign singleKey_145_raw = key_down[42];
  assign keyStatus_42_valid = singleKey_145_filtered_valid;
  assign keyStatus_42_payload = singleKey_145_filtered_payload;
  assign singleKey_146_raw = key_down[43];
  assign keyStatus_43_valid = singleKey_146_filtered_valid;
  assign keyStatus_43_payload = singleKey_146_filtered_payload;
  assign singleKey_147_raw = key_down[44];
  assign keyStatus_44_valid = singleKey_147_filtered_valid;
  assign keyStatus_44_payload = singleKey_147_filtered_payload;
  assign singleKey_148_raw = key_down[45];
  assign keyStatus_45_valid = singleKey_148_filtered_valid;
  assign keyStatus_45_payload = singleKey_148_filtered_payload;
  assign singleKey_149_raw = key_down[46];
  assign keyStatus_46_valid = singleKey_149_filtered_valid;
  assign keyStatus_46_payload = singleKey_149_filtered_payload;
  assign singleKey_150_raw = key_down[47];
  assign keyStatus_47_valid = singleKey_150_filtered_valid;
  assign keyStatus_47_payload = singleKey_150_filtered_payload;
  assign singleKey_151_raw = key_down[48];
  assign keyStatus_48_valid = singleKey_151_filtered_valid;
  assign keyStatus_48_payload = singleKey_151_filtered_payload;
  assign singleKey_152_raw = key_down[49];
  assign keyStatus_49_valid = singleKey_152_filtered_valid;
  assign keyStatus_49_payload = singleKey_152_filtered_payload;
  assign singleKey_153_raw = key_down[50];
  assign keyStatus_50_valid = singleKey_153_filtered_valid;
  assign keyStatus_50_payload = singleKey_153_filtered_payload;
  assign singleKey_154_raw = key_down[51];
  assign keyStatus_51_valid = singleKey_154_filtered_valid;
  assign keyStatus_51_payload = singleKey_154_filtered_payload;
  assign singleKey_155_raw = key_down[52];
  assign keyStatus_52_valid = singleKey_155_filtered_valid;
  assign keyStatus_52_payload = singleKey_155_filtered_payload;
  assign singleKey_156_raw = key_down[53];
  assign keyStatus_53_valid = singleKey_156_filtered_valid;
  assign keyStatus_53_payload = singleKey_156_filtered_payload;
  assign singleKey_157_raw = key_down[54];
  assign keyStatus_54_valid = singleKey_157_filtered_valid;
  assign keyStatus_54_payload = singleKey_157_filtered_payload;
  assign singleKey_158_raw = key_down[55];
  assign keyStatus_55_valid = singleKey_158_filtered_valid;
  assign keyStatus_55_payload = singleKey_158_filtered_payload;
  assign singleKey_159_raw = key_down[56];
  assign keyStatus_56_valid = singleKey_159_filtered_valid;
  assign keyStatus_56_payload = singleKey_159_filtered_payload;
  assign singleKey_160_raw = key_down[57];
  assign keyStatus_57_valid = singleKey_160_filtered_valid;
  assign keyStatus_57_payload = singleKey_160_filtered_payload;
  assign singleKey_161_raw = key_down[58];
  assign keyStatus_58_valid = singleKey_161_filtered_valid;
  assign keyStatus_58_payload = singleKey_161_filtered_payload;
  assign singleKey_162_raw = key_down[59];
  assign keyStatus_59_valid = singleKey_162_filtered_valid;
  assign keyStatus_59_payload = singleKey_162_filtered_payload;
  assign singleKey_163_raw = key_down[60];
  assign keyStatus_60_valid = singleKey_163_filtered_valid;
  assign keyStatus_60_payload = singleKey_163_filtered_payload;
  assign singleKey_164_raw = key_down[61];
  assign keyStatus_61_valid = singleKey_164_filtered_valid;
  assign keyStatus_61_payload = singleKey_164_filtered_payload;
  assign singleKey_165_raw = key_down[62];
  assign keyStatus_62_valid = singleKey_165_filtered_valid;
  assign keyStatus_62_payload = singleKey_165_filtered_payload;
  assign singleKey_166_raw = key_down[63];
  assign keyStatus_63_valid = singleKey_166_filtered_valid;
  assign keyStatus_63_payload = singleKey_166_filtered_payload;
  assign singleKey_167_raw = key_down[64];
  assign keyStatus_64_valid = singleKey_167_filtered_valid;
  assign keyStatus_64_payload = singleKey_167_filtered_payload;
  assign singleKey_168_raw = key_down[65];
  assign keyStatus_65_valid = singleKey_168_filtered_valid;
  assign keyStatus_65_payload = singleKey_168_filtered_payload;
  assign singleKey_169_raw = key_down[66];
  assign keyStatus_66_valid = singleKey_169_filtered_valid;
  assign keyStatus_66_payload = singleKey_169_filtered_payload;
  assign singleKey_170_raw = key_down[67];
  assign keyStatus_67_valid = singleKey_170_filtered_valid;
  assign keyStatus_67_payload = singleKey_170_filtered_payload;
  assign singleKey_171_raw = key_down[68];
  assign keyStatus_68_valid = singleKey_171_filtered_valid;
  assign keyStatus_68_payload = singleKey_171_filtered_payload;
  assign singleKey_172_raw = key_down[69];
  assign keyStatus_69_valid = singleKey_172_filtered_valid;
  assign keyStatus_69_payload = singleKey_172_filtered_payload;
  assign singleKey_173_raw = key_down[70];
  assign keyStatus_70_valid = singleKey_173_filtered_valid;
  assign keyStatus_70_payload = singleKey_173_filtered_payload;
  assign singleKey_174_raw = key_down[71];
  assign keyStatus_71_valid = singleKey_174_filtered_valid;
  assign keyStatus_71_payload = singleKey_174_filtered_payload;
  assign singleKey_175_raw = key_down[72];
  assign keyStatus_72_valid = singleKey_175_filtered_valid;
  assign keyStatus_72_payload = singleKey_175_filtered_payload;
  assign singleKey_176_raw = key_down[73];
  assign keyStatus_73_valid = singleKey_176_filtered_valid;
  assign keyStatus_73_payload = singleKey_176_filtered_payload;
  assign singleKey_177_raw = key_down[74];
  assign keyStatus_74_valid = singleKey_177_filtered_valid;
  assign keyStatus_74_payload = singleKey_177_filtered_payload;
  assign singleKey_178_raw = key_down[75];
  assign keyStatus_75_valid = singleKey_178_filtered_valid;
  assign keyStatus_75_payload = singleKey_178_filtered_payload;
  assign singleKey_179_raw = key_down[76];
  assign keyStatus_76_valid = singleKey_179_filtered_valid;
  assign keyStatus_76_payload = singleKey_179_filtered_payload;
  assign singleKey_180_raw = key_down[77];
  assign keyStatus_77_valid = singleKey_180_filtered_valid;
  assign keyStatus_77_payload = singleKey_180_filtered_payload;
  assign singleKey_181_raw = key_down[78];
  assign keyStatus_78_valid = singleKey_181_filtered_valid;
  assign keyStatus_78_payload = singleKey_181_filtered_payload;
  assign singleKey_182_raw = key_down[79];
  assign keyStatus_79_valid = singleKey_182_filtered_valid;
  assign keyStatus_79_payload = singleKey_182_filtered_payload;
  assign singleKey_183_raw = key_down[80];
  assign keyStatus_80_valid = singleKey_183_filtered_valid;
  assign keyStatus_80_payload = singleKey_183_filtered_payload;
  assign singleKey_184_raw = key_down[81];
  assign keyStatus_81_valid = singleKey_184_filtered_valid;
  assign keyStatus_81_payload = singleKey_184_filtered_payload;
  assign singleKey_185_raw = key_down[82];
  assign keyStatus_82_valid = singleKey_185_filtered_valid;
  assign keyStatus_82_payload = singleKey_185_filtered_payload;
  assign singleKey_186_raw = key_down[83];
  assign keyStatus_83_valid = singleKey_186_filtered_valid;
  assign keyStatus_83_payload = singleKey_186_filtered_payload;
  assign singleKey_187_raw = key_down[84];
  assign keyStatus_84_valid = singleKey_187_filtered_valid;
  assign keyStatus_84_payload = singleKey_187_filtered_payload;
  assign singleKey_188_raw = key_down[85];
  assign keyStatus_85_valid = singleKey_188_filtered_valid;
  assign keyStatus_85_payload = singleKey_188_filtered_payload;
  assign singleKey_189_raw = key_down[86];
  assign keyStatus_86_valid = singleKey_189_filtered_valid;
  assign keyStatus_86_payload = singleKey_189_filtered_payload;
  assign singleKey_190_raw = key_down[87];
  assign keyStatus_87_valid = singleKey_190_filtered_valid;
  assign keyStatus_87_payload = singleKey_190_filtered_payload;
  assign singleKey_191_raw = key_down[88];
  assign keyStatus_88_valid = singleKey_191_filtered_valid;
  assign keyStatus_88_payload = singleKey_191_filtered_payload;
  assign singleKey_192_raw = key_down[89];
  assign keyStatus_89_valid = singleKey_192_filtered_valid;
  assign keyStatus_89_payload = singleKey_192_filtered_payload;
  assign singleKey_193_raw = key_down[90];
  assign keyStatus_90_valid = singleKey_193_filtered_valid;
  assign keyStatus_90_payload = singleKey_193_filtered_payload;
  assign singleKey_194_raw = key_down[91];
  assign keyStatus_91_valid = singleKey_194_filtered_valid;
  assign keyStatus_91_payload = singleKey_194_filtered_payload;
  assign singleKey_195_raw = key_down[92];
  assign keyStatus_92_valid = singleKey_195_filtered_valid;
  assign keyStatus_92_payload = singleKey_195_filtered_payload;
  assign singleKey_196_raw = key_down[93];
  assign keyStatus_93_valid = singleKey_196_filtered_valid;
  assign keyStatus_93_payload = singleKey_196_filtered_payload;
  assign singleKey_197_raw = key_down[94];
  assign keyStatus_94_valid = singleKey_197_filtered_valid;
  assign keyStatus_94_payload = singleKey_197_filtered_payload;
  assign singleKey_198_raw = key_down[95];
  assign keyStatus_95_valid = singleKey_198_filtered_valid;
  assign keyStatus_95_payload = singleKey_198_filtered_payload;
  assign singleKey_199_raw = key_down[96];
  assign keyStatus_96_valid = singleKey_199_filtered_valid;
  assign keyStatus_96_payload = singleKey_199_filtered_payload;
  assign singleKey_200_raw = key_down[97];
  assign keyStatus_97_valid = singleKey_200_filtered_valid;
  assign keyStatus_97_payload = singleKey_200_filtered_payload;
  assign singleKey_201_raw = key_down[98];
  assign keyStatus_98_valid = singleKey_201_filtered_valid;
  assign keyStatus_98_payload = singleKey_201_filtered_payload;
  assign singleKey_202_raw = key_down[99];
  assign keyStatus_99_valid = singleKey_202_filtered_valid;
  assign keyStatus_99_payload = singleKey_202_filtered_payload;
  assign singleKey_203_raw = key_down[100];
  assign keyStatus_100_valid = singleKey_203_filtered_valid;
  assign keyStatus_100_payload = singleKey_203_filtered_payload;
  assign singleKey_204_raw = key_down[101];
  assign keyStatus_101_valid = singleKey_204_filtered_valid;
  assign keyStatus_101_payload = singleKey_204_filtered_payload;
  assign singleKey_205_raw = key_down[102];
  assign keyStatus_102_valid = singleKey_205_filtered_valid;
  assign keyStatus_102_payload = singleKey_205_filtered_payload;
  always @(posedge CLK_50 or posedge _zz_LED_R6) begin
    if(_zz_LED_R6) begin
      _zz_when_ClockDomain_l369 <= 15'h0;
      when_ClockDomain_l369_regNext <= 1'b0;
    end else begin
      _zz_when_ClockDomain_l369 <= (_zz_when_ClockDomain_l369 + 15'h0001);
      if(when_ClockDomain_l369) begin
        _zz_when_ClockDomain_l369 <= 15'h0;
      end
      when_ClockDomain_l369_regNext <= when_ClockDomain_l369;
    end
  end


endmodule

module UartCtrlRx_1 (
  input      [2:0]    io_configFrame_dataLength,
  input      [0:0]    io_configFrame_stop,
  input      [1:0]    io_configFrame_parity,
  input               io_samplingTick,
  output              io_read_valid,
  input               io_read_ready,
  output     [7:0]    io_read_payload,
  input               io_rxd,
  output              io_rts,
  output reg          io_error,
  output              io_break,
  input               CLK_50,
  input               _zz_LED_R6
);
  localparam UartStopType_ONE = 1'd0;
  localparam UartStopType_TWO = 1'd1;
  localparam UartParityType_NONE = 2'd0;
  localparam UartParityType_EVEN = 2'd1;
  localparam UartParityType_ODD = 2'd2;
  localparam UartCtrlRxState_IDLE = 3'd0;
  localparam UartCtrlRxState_START = 3'd1;
  localparam UartCtrlRxState_DATA = 3'd2;
  localparam UartCtrlRxState_PARITY = 3'd3;
  localparam UartCtrlRxState_STOP = 3'd4;

  wire                io_rxd_buffercc_io_dataOut;
  wire                _zz_sampler_value;
  wire                _zz_sampler_value_1;
  wire                _zz_sampler_value_2;
  wire                _zz_sampler_value_3;
  wire                _zz_sampler_value_4;
  wire                _zz_sampler_value_5;
  wire                _zz_sampler_value_6;
  wire       [2:0]    _zz_when_UartCtrlRx_l139;
  wire       [0:0]    _zz_when_UartCtrlRx_l139_1;
  reg                 _zz_io_rts;
  wire                sampler_synchroniser;
  wire                sampler_samples_0;
  reg                 sampler_samples_1;
  reg                 sampler_samples_2;
  reg                 sampler_samples_3;
  reg                 sampler_samples_4;
  reg                 sampler_value;
  reg                 sampler_tick;
  reg        [2:0]    bitTimer_counter;
  reg                 bitTimer_tick;
  wire                when_UartCtrlRx_l43;
  reg        [2:0]    bitCounter_value;
  reg        [6:0]    break_counter;
  wire                break_valid;
  wire                when_UartCtrlRx_l69;
  reg        [2:0]    stateMachine_state;
  reg                 stateMachine_parity;
  reg        [7:0]    stateMachine_shifter;
  reg                 stateMachine_validReg;
  wire                when_UartCtrlRx_l93;
  wire                when_UartCtrlRx_l103;
  wire                when_UartCtrlRx_l111;
  wire                when_UartCtrlRx_l113;
  wire                when_UartCtrlRx_l125;
  wire                when_UartCtrlRx_l136;
  wire                when_UartCtrlRx_l139;
  `ifndef SYNTHESIS
  reg [23:0] io_configFrame_stop_string;
  reg [31:0] io_configFrame_parity_string;
  reg [47:0] stateMachine_state_string;
  `endif


  assign _zz_when_UartCtrlRx_l139_1 = ((io_configFrame_stop == UartStopType_ONE) ? 1'b0 : 1'b1);
  assign _zz_when_UartCtrlRx_l139 = {2'd0, _zz_when_UartCtrlRx_l139_1};
  assign _zz_sampler_value = ((((1'b0 || ((_zz_sampler_value_1 && sampler_samples_1) && sampler_samples_2)) || (((_zz_sampler_value_2 && sampler_samples_0) && sampler_samples_1) && sampler_samples_3)) || (((1'b1 && sampler_samples_0) && sampler_samples_2) && sampler_samples_3)) || (((1'b1 && sampler_samples_1) && sampler_samples_2) && sampler_samples_3));
  assign _zz_sampler_value_3 = (((1'b1 && sampler_samples_0) && sampler_samples_1) && sampler_samples_4);
  assign _zz_sampler_value_4 = ((1'b1 && sampler_samples_0) && sampler_samples_2);
  assign _zz_sampler_value_5 = (1'b1 && sampler_samples_1);
  assign _zz_sampler_value_6 = 1'b1;
  assign _zz_sampler_value_1 = (1'b1 && sampler_samples_0);
  assign _zz_sampler_value_2 = 1'b1;
  BufferCC_2 io_rxd_buffercc (
    .io_dataIn  (io_rxd                    ), //i
    .io_dataOut (io_rxd_buffercc_io_dataOut), //o
    .CLK_50     (CLK_50                    ), //i
    ._zz_LED_R6 (_zz_LED_R6                )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_configFrame_stop)
      UartStopType_ONE : io_configFrame_stop_string = "ONE";
      UartStopType_TWO : io_configFrame_stop_string = "TWO";
      default : io_configFrame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_configFrame_parity)
      UartParityType_NONE : io_configFrame_parity_string = "NONE";
      UartParityType_EVEN : io_configFrame_parity_string = "EVEN";
      UartParityType_ODD : io_configFrame_parity_string = "ODD ";
      default : io_configFrame_parity_string = "????";
    endcase
  end
  always @(*) begin
    case(stateMachine_state)
      UartCtrlRxState_IDLE : stateMachine_state_string = "IDLE  ";
      UartCtrlRxState_START : stateMachine_state_string = "START ";
      UartCtrlRxState_DATA : stateMachine_state_string = "DATA  ";
      UartCtrlRxState_PARITY : stateMachine_state_string = "PARITY";
      UartCtrlRxState_STOP : stateMachine_state_string = "STOP  ";
      default : stateMachine_state_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    io_error = 1'b0;
    case(stateMachine_state)
      UartCtrlRxState_IDLE : begin
      end
      UartCtrlRxState_START : begin
      end
      UartCtrlRxState_DATA : begin
      end
      UartCtrlRxState_PARITY : begin
        if(bitTimer_tick) begin
          if(!when_UartCtrlRx_l125) begin
            io_error = 1'b1;
          end
        end
      end
      default : begin
        if(bitTimer_tick) begin
          if(when_UartCtrlRx_l136) begin
            io_error = 1'b1;
          end
        end
      end
    endcase
  end

  assign io_rts = _zz_io_rts;
  assign sampler_synchroniser = io_rxd_buffercc_io_dataOut;
  assign sampler_samples_0 = sampler_synchroniser;
  always @(*) begin
    bitTimer_tick = 1'b0;
    if(sampler_tick) begin
      if(when_UartCtrlRx_l43) begin
        bitTimer_tick = 1'b1;
      end
    end
  end

  assign when_UartCtrlRx_l43 = (bitTimer_counter == 3'b000);
  assign break_valid = (break_counter == 7'h68);
  assign when_UartCtrlRx_l69 = (io_samplingTick && (! break_valid));
  assign io_break = break_valid;
  assign io_read_valid = stateMachine_validReg;
  assign when_UartCtrlRx_l93 = ((sampler_tick && (! sampler_value)) && (! break_valid));
  assign when_UartCtrlRx_l103 = (sampler_value == 1'b1);
  assign when_UartCtrlRx_l111 = (bitCounter_value == io_configFrame_dataLength);
  assign when_UartCtrlRx_l113 = (io_configFrame_parity == UartParityType_NONE);
  assign when_UartCtrlRx_l125 = (stateMachine_parity == sampler_value);
  assign when_UartCtrlRx_l136 = (! sampler_value);
  assign when_UartCtrlRx_l139 = (bitCounter_value == _zz_when_UartCtrlRx_l139);
  assign io_read_payload = stateMachine_shifter;
  always @(posedge CLK_50 or posedge _zz_LED_R6) begin
    if(_zz_LED_R6) begin
      _zz_io_rts <= 1'b0;
      sampler_samples_1 <= 1'b1;
      sampler_samples_2 <= 1'b1;
      sampler_samples_3 <= 1'b1;
      sampler_samples_4 <= 1'b1;
      sampler_value <= 1'b1;
      sampler_tick <= 1'b0;
      break_counter <= 7'h0;
      stateMachine_state <= UartCtrlRxState_IDLE;
      stateMachine_validReg <= 1'b0;
    end else begin
      _zz_io_rts <= (! io_read_ready);
      if(io_samplingTick) begin
        sampler_samples_1 <= sampler_samples_0;
      end
      if(io_samplingTick) begin
        sampler_samples_2 <= sampler_samples_1;
      end
      if(io_samplingTick) begin
        sampler_samples_3 <= sampler_samples_2;
      end
      if(io_samplingTick) begin
        sampler_samples_4 <= sampler_samples_3;
      end
      sampler_value <= ((((((_zz_sampler_value || _zz_sampler_value_3) || (_zz_sampler_value_4 && sampler_samples_4)) || ((_zz_sampler_value_5 && sampler_samples_2) && sampler_samples_4)) || (((_zz_sampler_value_6 && sampler_samples_0) && sampler_samples_3) && sampler_samples_4)) || (((1'b1 && sampler_samples_1) && sampler_samples_3) && sampler_samples_4)) || (((1'b1 && sampler_samples_2) && sampler_samples_3) && sampler_samples_4));
      sampler_tick <= io_samplingTick;
      if(sampler_value) begin
        break_counter <= 7'h0;
      end else begin
        if(when_UartCtrlRx_l69) begin
          break_counter <= (break_counter + 7'h01);
        end
      end
      stateMachine_validReg <= 1'b0;
      case(stateMachine_state)
        UartCtrlRxState_IDLE : begin
          if(when_UartCtrlRx_l93) begin
            stateMachine_state <= UartCtrlRxState_START;
          end
        end
        UartCtrlRxState_START : begin
          if(bitTimer_tick) begin
            stateMachine_state <= UartCtrlRxState_DATA;
            if(when_UartCtrlRx_l103) begin
              stateMachine_state <= UartCtrlRxState_IDLE;
            end
          end
        end
        UartCtrlRxState_DATA : begin
          if(bitTimer_tick) begin
            if(when_UartCtrlRx_l111) begin
              if(when_UartCtrlRx_l113) begin
                stateMachine_state <= UartCtrlRxState_STOP;
                stateMachine_validReg <= 1'b1;
              end else begin
                stateMachine_state <= UartCtrlRxState_PARITY;
              end
            end
          end
        end
        UartCtrlRxState_PARITY : begin
          if(bitTimer_tick) begin
            if(when_UartCtrlRx_l125) begin
              stateMachine_state <= UartCtrlRxState_STOP;
              stateMachine_validReg <= 1'b1;
            end else begin
              stateMachine_state <= UartCtrlRxState_IDLE;
            end
          end
        end
        default : begin
          if(bitTimer_tick) begin
            if(when_UartCtrlRx_l136) begin
              stateMachine_state <= UartCtrlRxState_IDLE;
            end else begin
              if(when_UartCtrlRx_l139) begin
                stateMachine_state <= UartCtrlRxState_IDLE;
              end
            end
          end
        end
      endcase
    end
  end

  always @(posedge CLK_50) begin
    if(sampler_tick) begin
      bitTimer_counter <= (bitTimer_counter - 3'b001);
    end
    if(bitTimer_tick) begin
      bitCounter_value <= (bitCounter_value + 3'b001);
    end
    if(bitTimer_tick) begin
      stateMachine_parity <= (stateMachine_parity ^ sampler_value);
    end
    case(stateMachine_state)
      UartCtrlRxState_IDLE : begin
        if(when_UartCtrlRx_l93) begin
          bitTimer_counter <= 3'b010;
        end
      end
      UartCtrlRxState_START : begin
        if(bitTimer_tick) begin
          bitCounter_value <= 3'b000;
          stateMachine_parity <= (io_configFrame_parity == UartParityType_ODD);
        end
      end
      UartCtrlRxState_DATA : begin
        if(bitTimer_tick) begin
          stateMachine_shifter[bitCounter_value] <= sampler_value;
          if(when_UartCtrlRx_l111) begin
            bitCounter_value <= 3'b000;
          end
        end
      end
      UartCtrlRxState_PARITY : begin
        if(bitTimer_tick) begin
          bitCounter_value <= 3'b000;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module UartCtrlTx_1 (
  input      [2:0]    io_configFrame_dataLength,
  input      [0:0]    io_configFrame_stop,
  input      [1:0]    io_configFrame_parity,
  input               io_samplingTick,
  input               io_write_valid,
  output reg          io_write_ready,
  input      [7:0]    io_write_payload,
  input               io_cts,
  output              io_txd,
  input               io_break,
  input               CLK_50,
  input               _zz_LED_R6
);
  localparam UartStopType_ONE = 1'd0;
  localparam UartStopType_TWO = 1'd1;
  localparam UartParityType_NONE = 2'd0;
  localparam UartParityType_EVEN = 2'd1;
  localparam UartParityType_ODD = 2'd2;
  localparam UartCtrlTxState_IDLE = 3'd0;
  localparam UartCtrlTxState_START = 3'd1;
  localparam UartCtrlTxState_DATA = 3'd2;
  localparam UartCtrlTxState_PARITY = 3'd3;
  localparam UartCtrlTxState_STOP = 3'd4;

  wire       [2:0]    _zz_clockDivider_counter_valueNext;
  wire       [0:0]    _zz_clockDivider_counter_valueNext_1;
  wire       [2:0]    _zz_when_UartCtrlTx_l93;
  wire       [0:0]    _zz_when_UartCtrlTx_l93_1;
  reg                 clockDivider_counter_willIncrement;
  wire                clockDivider_counter_willClear;
  reg        [2:0]    clockDivider_counter_valueNext;
  reg        [2:0]    clockDivider_counter_value;
  wire                clockDivider_counter_willOverflowIfInc;
  wire                clockDivider_counter_willOverflow;
  reg        [2:0]    tickCounter_value;
  reg        [2:0]    stateMachine_state;
  reg                 stateMachine_parity;
  reg                 stateMachine_txd;
  wire                when_UartCtrlTx_l58;
  wire                when_UartCtrlTx_l73;
  wire                when_UartCtrlTx_l76;
  wire                when_UartCtrlTx_l93;
  wire       [2:0]    _zz_stateMachine_state;
  reg                 _zz_io_txd;
  `ifndef SYNTHESIS
  reg [23:0] io_configFrame_stop_string;
  reg [31:0] io_configFrame_parity_string;
  reg [47:0] stateMachine_state_string;
  reg [47:0] _zz_stateMachine_state_string;
  `endif


  assign _zz_clockDivider_counter_valueNext_1 = clockDivider_counter_willIncrement;
  assign _zz_clockDivider_counter_valueNext = {2'd0, _zz_clockDivider_counter_valueNext_1};
  assign _zz_when_UartCtrlTx_l93_1 = ((io_configFrame_stop == UartStopType_ONE) ? 1'b0 : 1'b1);
  assign _zz_when_UartCtrlTx_l93 = {2'd0, _zz_when_UartCtrlTx_l93_1};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_configFrame_stop)
      UartStopType_ONE : io_configFrame_stop_string = "ONE";
      UartStopType_TWO : io_configFrame_stop_string = "TWO";
      default : io_configFrame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_configFrame_parity)
      UartParityType_NONE : io_configFrame_parity_string = "NONE";
      UartParityType_EVEN : io_configFrame_parity_string = "EVEN";
      UartParityType_ODD : io_configFrame_parity_string = "ODD ";
      default : io_configFrame_parity_string = "????";
    endcase
  end
  always @(*) begin
    case(stateMachine_state)
      UartCtrlTxState_IDLE : stateMachine_state_string = "IDLE  ";
      UartCtrlTxState_START : stateMachine_state_string = "START ";
      UartCtrlTxState_DATA : stateMachine_state_string = "DATA  ";
      UartCtrlTxState_PARITY : stateMachine_state_string = "PARITY";
      UartCtrlTxState_STOP : stateMachine_state_string = "STOP  ";
      default : stateMachine_state_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_stateMachine_state)
      UartCtrlTxState_IDLE : _zz_stateMachine_state_string = "IDLE  ";
      UartCtrlTxState_START : _zz_stateMachine_state_string = "START ";
      UartCtrlTxState_DATA : _zz_stateMachine_state_string = "DATA  ";
      UartCtrlTxState_PARITY : _zz_stateMachine_state_string = "PARITY";
      UartCtrlTxState_STOP : _zz_stateMachine_state_string = "STOP  ";
      default : _zz_stateMachine_state_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    clockDivider_counter_willIncrement = 1'b0;
    if(io_samplingTick) begin
      clockDivider_counter_willIncrement = 1'b1;
    end
  end

  assign clockDivider_counter_willClear = 1'b0;
  assign clockDivider_counter_willOverflowIfInc = (clockDivider_counter_value == 3'b111);
  assign clockDivider_counter_willOverflow = (clockDivider_counter_willOverflowIfInc && clockDivider_counter_willIncrement);
  always @(*) begin
    clockDivider_counter_valueNext = (clockDivider_counter_value + _zz_clockDivider_counter_valueNext);
    if(clockDivider_counter_willClear) begin
      clockDivider_counter_valueNext = 3'b000;
    end
  end

  always @(*) begin
    stateMachine_txd = 1'b1;
    case(stateMachine_state)
      UartCtrlTxState_IDLE : begin
      end
      UartCtrlTxState_START : begin
        stateMachine_txd = 1'b0;
      end
      UartCtrlTxState_DATA : begin
        stateMachine_txd = io_write_payload[tickCounter_value];
      end
      UartCtrlTxState_PARITY : begin
        stateMachine_txd = stateMachine_parity;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_write_ready = io_break;
    case(stateMachine_state)
      UartCtrlTxState_IDLE : begin
      end
      UartCtrlTxState_START : begin
      end
      UartCtrlTxState_DATA : begin
        if(clockDivider_counter_willOverflow) begin
          if(when_UartCtrlTx_l73) begin
            io_write_ready = 1'b1;
          end
        end
      end
      UartCtrlTxState_PARITY : begin
      end
      default : begin
      end
    endcase
  end

  assign when_UartCtrlTx_l58 = ((io_write_valid && (! io_cts)) && clockDivider_counter_willOverflow);
  assign when_UartCtrlTx_l73 = (tickCounter_value == io_configFrame_dataLength);
  assign when_UartCtrlTx_l76 = (io_configFrame_parity == UartParityType_NONE);
  assign when_UartCtrlTx_l93 = (tickCounter_value == _zz_when_UartCtrlTx_l93);
  assign _zz_stateMachine_state = (io_write_valid ? UartCtrlTxState_START : UartCtrlTxState_IDLE);
  assign io_txd = _zz_io_txd;
  always @(posedge CLK_50 or posedge _zz_LED_R6) begin
    if(_zz_LED_R6) begin
      clockDivider_counter_value <= 3'b000;
      stateMachine_state <= UartCtrlTxState_IDLE;
      _zz_io_txd <= 1'b1;
    end else begin
      clockDivider_counter_value <= clockDivider_counter_valueNext;
      case(stateMachine_state)
        UartCtrlTxState_IDLE : begin
          if(when_UartCtrlTx_l58) begin
            stateMachine_state <= UartCtrlTxState_START;
          end
        end
        UartCtrlTxState_START : begin
          if(clockDivider_counter_willOverflow) begin
            stateMachine_state <= UartCtrlTxState_DATA;
          end
        end
        UartCtrlTxState_DATA : begin
          if(clockDivider_counter_willOverflow) begin
            if(when_UartCtrlTx_l73) begin
              if(when_UartCtrlTx_l76) begin
                stateMachine_state <= UartCtrlTxState_STOP;
              end else begin
                stateMachine_state <= UartCtrlTxState_PARITY;
              end
            end
          end
        end
        UartCtrlTxState_PARITY : begin
          if(clockDivider_counter_willOverflow) begin
            stateMachine_state <= UartCtrlTxState_STOP;
          end
        end
        default : begin
          if(clockDivider_counter_willOverflow) begin
            if(when_UartCtrlTx_l93) begin
              stateMachine_state <= _zz_stateMachine_state;
            end
          end
        end
      endcase
      _zz_io_txd <= (stateMachine_txd && (! io_break));
    end
  end

  always @(posedge CLK_50) begin
    if(clockDivider_counter_willOverflow) begin
      tickCounter_value <= (tickCounter_value + 3'b001);
    end
    if(clockDivider_counter_willOverflow) begin
      stateMachine_parity <= (stateMachine_parity ^ stateMachine_txd);
    end
    case(stateMachine_state)
      UartCtrlTxState_IDLE : begin
      end
      UartCtrlTxState_START : begin
        if(clockDivider_counter_willOverflow) begin
          stateMachine_parity <= (io_configFrame_parity == UartParityType_ODD);
          tickCounter_value <= 3'b000;
        end
      end
      UartCtrlTxState_DATA : begin
        if(clockDivider_counter_willOverflow) begin
          if(when_UartCtrlTx_l73) begin
            tickCounter_value <= 3'b000;
          end
        end
      end
      UartCtrlTxState_PARITY : begin
        if(clockDivider_counter_willOverflow) begin
          tickCounter_value <= 3'b000;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

//BufferCC_2 replaced by BufferCC_2

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

//SingleKey_102 replaced by SingleKey_102

module SingleKey_102 (
  input               raw,
  output              filtered_valid,
  output              filtered_payload,
  input               CLK_50,
  input               _zz_LED_R6,
  input               when_ClockDomain_l369_regNext
);

  reg        [1:0]    cnt;
  reg                 raw_regNext;
  wire                when_Debounce_l15;
  wire                when_Debounce_l16;
  reg                 _zz_filtered_valid;
  wire                when_Debounce_l18;
  reg                 _zz_filtered_payload;

  assign when_Debounce_l15 = (raw ^ raw_regNext);
  assign when_Debounce_l16 = (cnt != 2'b00);
  assign filtered_valid = _zz_filtered_valid;
  assign when_Debounce_l18 = (cnt == 2'b01);
  assign filtered_payload = _zz_filtered_payload;
  always @(posedge CLK_50 or posedge _zz_LED_R6) begin
    if(_zz_LED_R6) begin
      cnt <= 2'b11;
    end else begin
      if(when_ClockDomain_l369_regNext) begin
        if(when_Debounce_l15) begin
          cnt <= 2'b11;
        end
        if(when_Debounce_l16) begin
          cnt <= (cnt - 2'b01);
        end
      end
    end
  end

  always @(posedge CLK_50) begin
    if(when_ClockDomain_l369_regNext) begin
      raw_regNext <= raw;
      _zz_filtered_valid <= (cnt == 2'b01);
      if(when_Debounce_l18) begin
        _zz_filtered_payload <= (! raw);
      end
    end
  end


endmodule

module BufferCC_2 (
  input               io_dataIn,
  output              io_dataOut,
  input               CLK_50,
  input               _zz_LED_R6
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge CLK_50 or posedge _zz_LED_R6) begin
    if(_zz_LED_R6) begin
      buffers_0 <= 1'b0;
      buffers_1 <= 1'b0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule
