// Generator : SpinalHDL v1.8.0b    git head : 761a30e521263983ddf14de3592f7a9f38bf0589
// Component : top4
// Git hash  : aa75c98d3aae6e7fc40f8bd4693eb03b16e38926

`timescale 1ns/1ps

module top4 (
  input               io_a,
  output              io_b
);


  assign io_b = io_a;

endmodule
