// Generator : SpinalHDL v1.8.0b    git head : 761a30e521263983ddf14de3592f7a9f38bf0589
// Component : MyTry
// Git hash  : 83b5023813df2ca722096581cf13ad25bd8ea94d

`timescale 1ns/1ps

module MyTry (
  input               io_a,
  output              io_b
);


  assign io_b = io_a;

endmodule
